

.subckt TL_MS1 1 2 ngnd length=0.00643382


WTL1 1 ngnd 2 ngnd n=1 RLGCfile=G6Q3.rlc l='length'



.ends TL_MS1
