

.subckt TL_1 1 2 ngnd length=0.0020447


WTL1 1 ngnd 2 ngnd n=1 RLGCfile=w6l2.rlc l='length'



.ends TL_1
