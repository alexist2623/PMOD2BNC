********************************************************************************
*
* LTSPICE MODEL FOR IBIS MODEL(S)
* MODELING DATE: 20230619012917
* GENERAETD BY BPRO: http://www.spisim.com
*
* NOTE: ramp data in .ibs model is used in this converted spice model.
*       VT waveform based conversion will yield more accurate result.
*
********************************************************************************


******************************** BEGIN *****************************************
* ORIG. MDL: C:\Jeonghyun\GIT\PMOD2BNC\IBIS\spartan7_v1.3\spartan7\spartan7.ibs;LVCMOS33_S_8_HR;TYP
* TERMINALS: INPUT OUTPUT VCC VSS ENABLE

.SUBCKT LVCMOS33_S_8_HR_TYP NINP NOUT NVCC NVSS NENB

* POWER-ON SOURCE



* INPUT CONTROL
B1 N820 0 V= ((V(NINP) > 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0
B2 N830 0 V= ((V(NINP) < 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0

* RAMP RATE CONTROL
* RISERMP = 2.898695E5 = 1.0878/3.1532n
* FALLRMP = 1.001648E5 = 1.0920/1.0938n

B3 NVCC N850 I= (V(N830) > 0.5)? 0 : V(NVCC, N850) / 1.001648E5
B4 N840 NVSS I= (V(N820) > 0.5)? 0 : V(N840, NVSS) / 2.898695E5
C1 NVCC N850 1F
C2 N840 NVSS 1F
S1 N220 N850 0 N820 SMOD
S2 N840 N220 0 N830 SMOD

G1 N008 NVSS N002 N008 1
G2 NVCC N008 N008 N003 1
R1 N006 NVSS 1
R2 NVCC N006 1

* PU/PD/PC/GC BRANCH
XASRC_PD N002 NVSS N008 N840 LVCMOS33_S_8_HR_PULLDOWN_TYP
XASRC_PU N003 NVCC N850 N008 LVCMOS33_S_8_HR_PULLUP_TYP
XASRC_PC N006 NVCC NVCC N006 LVCMOS33_S_8_HR_POWER_CLAMP_TYP
XASRC_GC N006 NVSS N006 NVSS LVCMOS33_S_8_HR_GND_CLAMP_TYP

* PACKAGE PARASITICS:
ROPKG N001 NOUT 3.345000E-1
COPKG NOUT NVSS 7.200000E-13
LOPKG N005 N001 4.350000E-9
CCOMP N005 NVSS 5.230000E-12

* Voltage Sources for measuring currents
V5 N006 N005 0
V6 N008 N006 0
V7 N220 N008 0
.ENDS

* PU BRANCH
.SUBCKT LVCMOS33_S_8_HR_PULLUP_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -3.300000E0)? 2.867000E-2:
+ (V(1,2) < -3.200000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -3.100000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -3.000000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.900000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.800000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.700000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.600000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.500000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.400000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.300000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.200000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.100000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -2.000000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.900000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.800000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.700000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.600000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.500000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) + 2.867000E-2:
+ (V(1,2) < -8.000000E-1)? -2.370000E-2 * V(1,2) + 7.340000E-3:
+ (V(1,2) < -7.000000E-1)? -4.700000E-3 * V(1,2) + 2.254000E-2:
+ (V(1,2) < -6.000000E-1)? -1.420000E-2 * V(1,2) + 1.589000E-2:
+ (V(1,2) < -5.000000E-1)? -2.994000E-2 * V(1,2) + 6.446000E-3:
+ (V(1,2) < -4.000000E-1)? -1.504000E-2 * V(1,2) + 1.389600E-2:
+ (V(1,2) < -3.000000E-1)? -4.050300E-2 * V(1,2) + 3.710800E-3:
+ (V(1,2) < -2.000000E-1)? -5.671000E-2 * V(1,2) - 1.151300E-3:
+ (V(1,2) < -1.000000E-1)? -5.080900E-2 * V(1,2) + 2.890000E-5:
+ (V(1,2) < 0.000000E0)? -4.639500E-2 * V(1,2) + 4.703000E-4:
+ (V(1,2) < 1.000000E-1)? -4.422300E-2 * V(1,2) + 4.703000E-4:
+ (V(1,2) < 2.000000E-1)? -4.423000E-2 * V(1,2) + 4.710000E-4:
+ (V(1,2) < 3.000000E-1)? -4.425000E-2 * V(1,2) + 4.750000E-4:
+ (V(1,2) < 4.000000E-1)? -4.420000E-2 * V(1,2) + 4.600000E-4:
+ (V(1,2) < 5.000000E-1)? -3.320000E-2 * V(1,2) - 3.940000E-3:
+ (V(1,2) < 6.000000E-1)? -2.850000E-2 * V(1,2) - 6.290000E-3:
+ (V(1,2) < 7.000000E-1)? -2.850000E-2 * V(1,2) - 6.290000E-3:
+ (V(1,2) < 8.000000E-1)? -2.850000E-2 * V(1,2) - 6.290000E-3:
+ (V(1,2) < 9.000000E-1)? -1.940000E-2 * V(1,2) - 1.357000E-2:
+ (V(1,2) < 1.000000E0)? -1.640000E-2 * V(1,2) - 1.627000E-2:
+ (V(1,2) < 1.100000E0)? -1.560000E-2 * V(1,2) - 1.707000E-2:
+ (V(1,2) < 1.200000E0)? -8.800000E-3 * V(1,2) - 2.455000E-2:
+ (V(1,2) < 1.300000E0)? -6.700000E-3 * V(1,2) - 2.707000E-2:
+ (V(1,2) < 1.400000E0)? -3.700000E-3 * V(1,2) - 3.097000E-2:
+ (V(1,2) < 1.500000E0)? -2.400000E-3 * V(1,2) - 3.279000E-2:
+ (V(1,2) < 1.600000E0)? -2.000000E-3 * V(1,2) - 3.339000E-2:
+ (V(1,2) < 1.700000E0)? -1.600000E-3 * V(1,2) - 3.403000E-2:
+ (V(1,2) < 1.800000E0)? -1.300000E-3 * V(1,2) - 3.454000E-2:
+ (V(1,2) < 1.900000E0)? -1.300000E-3 * V(1,2) - 3.454000E-2:
+ (V(1,2) < 2.000000E0)? -1.100000E-3 * V(1,2) - 3.492000E-2:
+ (V(1,2) < 2.100000E0)? -1.100000E-3 * V(1,2) - 3.492000E-2:
+ (V(1,2) < 2.200000E0)? -1.000000E-3 * V(1,2) - 3.513000E-2:
+ (V(1,2) < 2.300000E0)? -9.000000E-4 * V(1,2) - 3.535000E-2:
+ (V(1,2) < 2.400000E0)? -5.720000E-2 * V(1,2) + 9.414000E-2:
+ (V(1,2) < 2.500000E0)? -6.000000E-4 * V(1,2) - 4.170000E-2:
+ (V(1,2) < 2.600000E0)? -6.000000E-4 * V(1,2) - 4.170000E-2:
+ (V(1,2) < 2.700000E0)? -6.000000E-4 * V(1,2) - 4.170000E-2:
+ (V(1,2) < 2.800000E0)? -5.000000E-4 * V(1,2) - 4.197000E-2:
+ (V(1,2) < 2.900000E0)? -5.000000E-4 * V(1,2) - 4.197000E-2:
+ (V(1,2) < 3.000000E0)? -5.000000E-4 * V(1,2) - 4.197000E-2:
+ (V(1,2) < 3.100000E0)? -6.000000E-4 * V(1,2) - 4.167000E-2:
+ (V(1,2) < 3.200000E0)? -4.000000E-4 * V(1,2) - 4.229000E-2:
+ (V(1,2) < 3.300000E0)? -5.000000E-4 * V(1,2) - 4.197000E-2:
+ (V(1,2) < 3.400000E0)? -4.990000E-4 * V(1,2) - 4.197330E-2:
+ (V(1,2) < 3.500000E0)? -4.870000E-4 * V(1,2) - 4.201410E-2:
+ (V(1,2) < 3.600000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 3.700000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 3.800000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 3.900000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.000000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.100000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.200000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.300000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.400000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.500000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.600000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.700000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.800000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 4.900000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.000000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.100000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.200000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.300000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.400000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.500000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.600000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.700000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.800000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 5.900000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 6.000000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 6.100000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 6.200000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 6.300000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 6.400000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 6.500000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ (V(1,2) < 6.600000E0)? -0.000000E0 * V(1,2) - 4.371860E-2:
+ -4.371860E-2 
.ENDS

* PD BRANCH
.SUBCKT LVCMOS33_S_8_HR_PULLDOWN_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -3.300000E0)? -2.644000E-2:
+ (V(1,2) < -3.200000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -3.100000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -3.000000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.900000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.800000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.700000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.600000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.500000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.400000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.300000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.200000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.100000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -2.000000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.900000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.800000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.700000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.600000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.500000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -8.000000E-1)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -7.000000E-1)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -6.000000E-1)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -5.000000E-1)? -0.000000E0 * V(1,2) - 2.644000E-2:
+ (V(1,2) < -4.000000E-1)? 4.466000E-3 * V(1,2) - 2.420700E-2:
+ (V(1,2) < -3.000000E-1)? 6.576300E-2 * V(1,2) + 3.118000E-4:
+ (V(1,2) < -2.000000E-1)? 6.586300E-2 * V(1,2) + 3.418000E-4:
+ (V(1,2) < -1.000000E-1)? 6.577300E-2 * V(1,2) + 3.238000E-4:
+ (V(1,2) < 0.000000E0)? 6.579500E-2 * V(1,2) + 3.260000E-4:
+ (V(1,2) < 1.000000E-1)? 6.595500E-2 * V(1,2) + 3.260000E-4:
+ (V(1,2) < 2.000000E-1)? 6.047700E-2 * V(1,2) + 8.738000E-4:
+ (V(1,2) < 3.000000E-1)? 5.250000E-2 * V(1,2) + 2.469200E-3:
+ (V(1,2) < 4.000000E-1)? 4.440000E-2 * V(1,2) + 4.899200E-3:
+ (V(1,2) < 5.000000E-1)? 3.650000E-2 * V(1,2) + 8.059200E-3:
+ (V(1,2) < 6.000000E-1)? 2.880000E-2 * V(1,2) + 1.190920E-2:
+ (V(1,2) < 7.000000E-1)? 2.360000E-2 * V(1,2) + 1.502920E-2:
+ (V(1,2) < 8.000000E-1)? 1.580000E-2 * V(1,2) + 2.048920E-2:
+ (V(1,2) < 9.000000E-1)? 1.490100E-2 * V(1,2) + 2.120840E-2:
+ (V(1,2) < 1.000000E0)? 7.500000E-3 * V(1,2) + 2.786930E-2:
+ (V(1,2) < 1.100000E0)? 4.700000E-3 * V(1,2) + 3.066930E-2:
+ (V(1,2) < 1.200000E0)? 2.700000E-3 * V(1,2) + 3.286930E-2:
+ (V(1,2) < 1.300000E0)? 1.800000E-3 * V(1,2) + 3.394930E-2:
+ (V(1,2) < 1.400000E0)? 1.301000E-3 * V(1,2) + 3.459800E-2:
+ (V(1,2) < 1.500000E0)? 6.000000E-4 * V(1,2) + 3.557940E-2:
+ (V(1,2) < 1.600000E0)? 6.000000E-4 * V(1,2) + 3.557940E-2:
+ (V(1,2) < 1.700000E0)? 4.000000E-4 * V(1,2) + 3.589940E-2:
+ (V(1,2) < 1.800000E0)? 4.000000E-4 * V(1,2) + 3.589940E-2:
+ (V(1,2) < 1.900000E0)? 4.000000E-4 * V(1,2) + 3.589940E-2:
+ (V(1,2) < 2.000000E0)? 3.000000E-4 * V(1,2) + 3.608940E-2:
+ (V(1,2) < 2.100000E0)? 2.990000E-4 * V(1,2) + 3.609140E-2:
+ (V(1,2) < 2.200000E0)? 4.000000E-4 * V(1,2) + 3.587930E-2:
+ (V(1,2) < 2.300000E0)? 2.740000E-2 * V(1,2) - 2.352070E-2:
+ (V(1,2) < 2.400000E0)? 3.000000E-4 * V(1,2) + 3.880930E-2:
+ (V(1,2) < 2.500000E0)? 2.990000E-4 * V(1,2) + 3.881170E-2:
+ (V(1,2) < 2.600000E0)? 2.000000E-4 * V(1,2) + 3.905920E-2:
+ (V(1,2) < 2.700000E0)? 3.000000E-4 * V(1,2) + 3.879920E-2:
+ (V(1,2) < 2.800000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 2.900000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.000000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.100000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.200000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.300000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.400000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.500000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.600000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.700000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.800000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 3.900000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.000000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.100000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.200000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.300000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.400000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.500000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.600000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.700000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.800000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 4.900000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.000000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.100000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.200000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.300000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.400000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.500000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.600000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.700000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.800000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 5.900000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 6.000000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 6.100000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 6.200000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 6.300000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 6.400000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 6.500000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ (V(1,2) < 6.600000E0)? -0.000000E0 * V(1,2) + 3.960920E-2:
+ 3.960920E-2 
.ENDS

* PC BRANCH
.SUBCKT LVCMOS33_S_8_HR_POWER_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -3.280000E0)? 3.564000E0:
+ (V(1,2) < -3.240000E0)? -1.550000E0 * V(1,2) - 1.520000E0:
+ (V(1,2) < -3.200000E0)? -1.525000E0 * V(1,2) - 1.439000E0:
+ (V(1,2) < -3.160000E0)? -1.550000E0 * V(1,2) - 1.519000E0:
+ (V(1,2) < -3.120000E0)? -1.525000E0 * V(1,2) - 1.440000E0:
+ (V(1,2) < -3.080000E0)? -1.550000E0 * V(1,2) - 1.518000E0:
+ (V(1,2) < -3.040000E0)? -1.525000E0 * V(1,2) - 1.441000E0:
+ (V(1,2) < -3.000000E0)? -1.550000E0 * V(1,2) - 1.517000E0:
+ (V(1,2) < -2.960000E0)? -1.525000E0 * V(1,2) - 1.442000E0:
+ (V(1,2) < -2.920000E0)? -1.550000E0 * V(1,2) - 1.516000E0:
+ (V(1,2) < -2.880000E0)? -1.525000E0 * V(1,2) - 1.443000E0:
+ (V(1,2) < -2.840000E0)? -1.550000E0 * V(1,2) - 1.515000E0:
+ (V(1,2) < -2.800000E0)? -1.525000E0 * V(1,2) - 1.444000E0:
+ (V(1,2) < -2.760000E0)? -1.525000E0 * V(1,2) - 1.444000E0:
+ (V(1,2) < -2.720000E0)? -1.550000E0 * V(1,2) - 1.513000E0:
+ (V(1,2) < -2.680000E0)? -1.525000E0 * V(1,2) - 1.445000E0:
+ (V(1,2) < -2.640000E0)? -1.550000E0 * V(1,2) - 1.512000E0:
+ (V(1,2) < -2.600000E0)? -1.525000E0 * V(1,2) - 1.446000E0:
+ (V(1,2) < -2.560000E0)? -1.550000E0 * V(1,2) - 1.511000E0:
+ (V(1,2) < -2.520000E0)? -1.525000E0 * V(1,2) - 1.447000E0:
+ (V(1,2) < -2.480000E0)? -1.550000E0 * V(1,2) - 1.510000E0:
+ (V(1,2) < -2.440000E0)? -1.525000E0 * V(1,2) - 1.448000E0:
+ (V(1,2) < -2.400000E0)? -1.550000E0 * V(1,2) - 1.509000E0:
+ (V(1,2) < -2.360000E0)? -1.525000E0 * V(1,2) - 1.449000E0:
+ (V(1,2) < -2.320000E0)? -1.550000E0 * V(1,2) - 1.508000E0:
+ (V(1,2) < -2.280000E0)? -1.525000E0 * V(1,2) - 1.450000E0:
+ (V(1,2) < -2.240000E0)? -1.525000E0 * V(1,2) - 1.450000E0:
+ (V(1,2) < -2.200000E0)? -1.550000E0 * V(1,2) - 1.506000E0:
+ (V(1,2) < -2.160000E0)? -1.525000E0 * V(1,2) - 1.451000E0:
+ (V(1,2) < -2.120000E0)? -1.550000E0 * V(1,2) - 1.505000E0:
+ (V(1,2) < -2.080000E0)? -1.525000E0 * V(1,2) - 1.452000E0:
+ (V(1,2) < -2.040000E0)? -1.550000E0 * V(1,2) - 1.504000E0:
+ (V(1,2) < -2.000000E0)? -1.525000E0 * V(1,2) - 1.453000E0:
+ (V(1,2) < -1.960000E0)? -1.550000E0 * V(1,2) - 1.503000E0:
+ (V(1,2) < -1.920000E0)? -1.525000E0 * V(1,2) - 1.454000E0:
+ (V(1,2) < -1.880000E0)? -1.550000E0 * V(1,2) - 1.502000E0:
+ (V(1,2) < -1.840000E0)? -1.525000E0 * V(1,2) - 1.455000E0:
+ (V(1,2) < -1.800000E0)? -1.525000E0 * V(1,2) - 1.455000E0:
+ (V(1,2) < -1.760000E0)? -1.550000E0 * V(1,2) - 1.500000E0:
+ (V(1,2) < -1.720000E0)? -1.525000E0 * V(1,2) - 1.456000E0:
+ (V(1,2) < -1.680000E0)? -1.550000E0 * V(1,2) - 1.499000E0:
+ (V(1,2) < -1.640000E0)? -1.525000E0 * V(1,2) - 1.457000E0:
+ (V(1,2) < -1.600000E0)? -1.532500E0 * V(1,2) - 1.469300E0:
+ (V(1,2) < -1.560000E0)? -1.535000E0 * V(1,2) - 1.473300E0:
+ (V(1,2) < -1.520000E0)? -1.532500E0 * V(1,2) - 1.469400E0:
+ (V(1,2) < -1.480000E0)? -1.532500E0 * V(1,2) - 1.469400E0:
+ (V(1,2) < -1.440000E0)? -1.530000E0 * V(1,2) - 1.465700E0:
+ (V(1,2) < -1.400000E0)? -1.530000E0 * V(1,2) - 1.465700E0:
+ (V(1,2) < -1.360000E0)? -1.532500E0 * V(1,2) - 1.469200E0:
+ (V(1,2) < -1.320000E0)? -1.495000E0 * V(1,2) - 1.418200E0:
+ (V(1,2) < -1.280000E0)? -1.462500E0 * V(1,2) - 1.375300E0:
+ (V(1,2) < -1.240000E0)? -1.462500E0 * V(1,2) - 1.375300E0:
+ (V(1,2) < -1.200000E0)? -1.465000E0 * V(1,2) - 1.378400E0:
+ (V(1,2) < -1.160000E0)? -1.462500E0 * V(1,2) - 1.375400E0:
+ (V(1,2) < -1.120000E0)? -1.370000E0 * V(1,2) - 1.268100E0:
+ (V(1,2) < -1.080000E0)? -1.290000E0 * V(1,2) - 1.178500E0:
+ (V(1,2) < -1.040000E0)? -1.292500E0 * V(1,2) - 1.181200E0:
+ (V(1,2) < -1.000000E0)? -1.125000E0 * V(1,2) - 1.007000E0:
+ (V(1,2) < -9.600000E-1)? -9.242500E-1 * V(1,2) - 8.062500E-1:
+ (V(1,2) < -9.200000E-1)? -6.375000E-1 * V(1,2) - 5.309700E-1:
+ (V(1,2) < -8.800000E-1)? -3.537500E-1 * V(1,2) - 2.699200E-1:
+ (V(1,2) < -8.400000E-1)? -2.055000E-1 * V(1,2) - 1.394600E-1:
+ (V(1,2) < -8.000000E-1)? -1.277500E-1 * V(1,2) - 7.415000E-2:
+ (V(1,2) < -7.600000E-1)? -8.875000E-2 * V(1,2) - 4.295000E-2:
+ (V(1,2) < -7.200000E-1)? -8.450000E-2 * V(1,2) - 3.972000E-2:
+ (V(1,2) < -6.800000E-1)? -8.425000E-2 * V(1,2) - 3.954000E-2:
+ (V(1,2) < -6.400000E-1)? -8.450000E-2 * V(1,2) - 3.971000E-2:
+ (V(1,2) < -6.000000E-1)? -8.450000E-2 * V(1,2) - 3.971000E-2:
+ (V(1,2) < -5.600000E-1)? -5.180000E-2 * V(1,2) - 2.009000E-2:
+ (V(1,2) < -5.200000E-1)? -4.835000E-2 * V(1,2) - 1.815800E-2:
+ (V(1,2) < -4.800000E-1)? -4.835000E-2 * V(1,2) - 1.815800E-2:
+ (V(1,2) < -4.400000E-1)? -4.832500E-2 * V(1,2) - 1.814600E-2:
+ (V(1,2) < -4.000000E-1)? -4.835000E-2 * V(1,2) - 1.815700E-2:
+ (V(1,2) < -3.600000E-1)? -1.004000E-2 * V(1,2) - 2.833000E-3:
+ (V(1,2) < -3.200000E-1)? -6.087500E-3 * V(1,2) - 1.410100E-3:
+ (V(1,2) < -2.800000E-1)? -6.087500E-3 * V(1,2) - 1.410100E-3:
+ (V(1,2) < -2.400000E-1)? -6.087000E-3 * V(1,2) - 1.409960E-3:
+ (V(1,2) < -2.000000E-1)? -1.121825E-3 * V(1,2) - 2.183180E-4:
+ (V(1,2) < -1.600000E-1)? -6.620000E-5 * V(1,2) - 7.193000E-6:
+ (V(1,2) < -1.200000E-1)? -6.618500E-5 * V(1,2) - 7.190600E-6:
+ (V(1,2) < -8.000000E-2)? -1.682575E-5 * V(1,2) - 1.267490E-6:
+ (V(1,2) < -4.000000E-2)? -1.230000E-6 * V(1,2) - 1.983000E-8:
+ (V(1,2) < 0.000000E0)? -2.442500E-7 * V(1,2) + 1.960000E-8:
+ 1.960000E-8 
.ENDS

* GC BRANCH
.SUBCKT LVCMOS33_S_8_HR_GND_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -3.300000E0)? -3.592000E0:
+ (V(1,2) < -3.230000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -3.160000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -3.090000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -3.020000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -2.950000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -2.880000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -2.810000E0)? 1.514286E0 * V(1,2) + 1.411143E0:
+ (V(1,2) < -2.740000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.670000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.600000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.530000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.460000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.390000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.320000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.250000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.180000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.110000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.040000E0)? 1.514286E0 * V(1,2) + 1.421143E0:
+ (V(1,2) < -1.970000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.900000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.830000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.760000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.690000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.620000E0)? 1.514286E0 * V(1,2) + 1.426143E0:
+ (V(1,2) < -1.550000E0)? 1.498571E0 * V(1,2) + 1.400686E0:
+ (V(1,2) < -1.480000E0)? 1.500000E0 * V(1,2) + 1.402900E0:
+ (V(1,2) < -1.410000E0)? 1.500000E0 * V(1,2) + 1.402900E0:
+ (V(1,2) < -1.340000E0)? 1.501429E0 * V(1,2) + 1.404914E0:
+ (V(1,2) < -1.270000E0)? 1.457143E0 * V(1,2) + 1.345571E0:
+ (V(1,2) < -1.200000E0)? 1.201429E0 * V(1,2) + 1.020814E0:
+ (V(1,2) < -1.130000E0)? 1.200000E0 * V(1,2) + 1.019100E0:
+ (V(1,2) < -1.060000E0)? 1.201429E0 * V(1,2) + 1.020714E0:
+ (V(1,2) < -9.900000E-1)? 1.200000E0 * V(1,2) + 1.019200E0:
+ (V(1,2) < -9.200000E-1)? 1.092857E0 * V(1,2) + 9.131286E-1:
+ (V(1,2) < -8.500000E-1)? 4.321429E-1 * V(1,2) + 3.052714E-1:
+ (V(1,2) < -7.800000E-1)? 2.414286E-1 * V(1,2) + 1.431643E-1:
+ (V(1,2) < -7.100000E-1)? 1.680000E-1 * V(1,2) + 8.589000E-2:
+ (V(1,2) < -6.400000E-1)? 1.680000E-1 * V(1,2) + 8.589000E-2:
+ (V(1,2) < -5.700000E-1)? 1.198571E-1 * V(1,2) + 5.507857E-2:
+ (V(1,2) < -5.000000E-1)? 9.605714E-2 * V(1,2) + 4.151257E-2:
+ (V(1,2) < -4.300000E-1)? 7.432857E-2 * V(1,2) + 3.064829E-2:
+ (V(1,2) < -3.600000E-1)? 1.553571E-2 * V(1,2) + 5.367357E-3:
+ (V(1,2) < -2.900000E-1)? 2.758286E-3 * V(1,2) + 7.674829E-4:
+ (V(1,2) < -2.200000E-1)? 3.637143E-4 * V(1,2) + 7.305714E-5:
+ (V(1,2) < -1.500000E-1)? 8.860714E-5 * V(1,2) + 1.253357E-5:
+ (V(1,2) < -8.000000E-2)? 1.035829E-5 * V(1,2) + 7.962429E-7:
+ (V(1,2) < -1.000000E-2)? 2.591429E-7 * V(1,2) - 1.168857E-8:
+ (V(1,2) < 6.000000E-2)? 2.914286E-8 * V(1,2) - 1.398857E-8:
+ (V(1,2) < 1.300000E-1)? 1.228571E-8 * V(1,2) - 1.297714E-8:
+ (V(1,2) < 2.000000E-1)? 9.000000E-9 * V(1,2) - 1.255000E-8:
+ (V(1,2) < 2.700000E-1)? 6.857143E-9 * V(1,2) - 1.212143E-8:
+ (V(1,2) < 3.400000E-1)? 6.342857E-9 * V(1,2) - 1.198257E-8:
+ (V(1,2) < 4.100000E-1)? 5.857143E-9 * V(1,2) - 1.181743E-8:
+ (V(1,2) < 4.800000E-1)? 5.842857E-9 * V(1,2) - 1.181157E-8:
+ (V(1,2) < 5.500000E-1)? 5.614286E-9 * V(1,2) - 1.170186E-8:
+ (V(1,2) < 6.200000E-1)? 5.557143E-9 * V(1,2) - 1.167043E-8:
+ (V(1,2) < 6.900000E-1)? 5.428571E-9 * V(1,2) - 1.159071E-8:
+ (V(1,2) < 7.600000E-1)? 5.414286E-9 * V(1,2) - 1.158086E-8:
+ (V(1,2) < 8.300000E-1)? 5.414286E-9 * V(1,2) - 1.158086E-8:
+ (V(1,2) < 9.000000E-1)? 5.400000E-9 * V(1,2) - 1.156900E-8:
+ (V(1,2) < 9.700000E-1)? 5.385714E-9 * V(1,2) - 1.155614E-8:
+ (V(1,2) < 1.040000E0)? 5.414286E-9 * V(1,2) - 1.158386E-8:
+ (V(1,2) < 1.110000E0)? 5.400000E-9 * V(1,2) - 1.156900E-8:
+ (V(1,2) < 1.180000E0)? 5.371429E-9 * V(1,2) - 1.153729E-8:
+ (V(1,2) < 1.250000E0)? 5.328571E-9 * V(1,2) - 1.148671E-8:
+ (V(1,2) < 1.320000E0)? 4.971429E-9 * V(1,2) - 1.104029E-8:
+ (V(1,2) < 1.390000E0)? 5.100000E-9 * V(1,2) - 1.121000E-8:
+ (V(1,2) < 1.460000E0)? 5.457143E-9 * V(1,2) - 1.170643E-8:
+ (V(1,2) < 1.530000E0)? 7.528571E-9 * V(1,2) - 1.473071E-8:
+ (V(1,2) < 1.600000E0)? 9.871429E-9 * V(1,2) - 1.831529E-8:
+ (V(1,2) < 1.670000E0)? 1.102857E-8 * V(1,2) - 2.016671E-8:
+ (V(1,2) < 1.740000E0)? 1.127143E-8 * V(1,2) - 2.057229E-8:
+ (V(1,2) < 1.810000E0)? 9.470000E-9 * V(1,2) - 1.743780E-8:
+ (V(1,2) < 1.880000E0)? 1.198429E-8 * V(1,2) - 2.198866E-8:
+ (V(1,2) < 1.950000E0)? 1.454571E-8 * V(1,2) - 2.680414E-8:
+ (V(1,2) < 2.020000E0)? 7.100000E-9 * V(1,2) - 1.228500E-8:
+ (V(1,2) < 2.090000E0)? 7.900000E-9 * V(1,2) - 1.390100E-8:
+ (V(1,2) < 2.160000E0)? 8.057143E-9 * V(1,2) - 1.422943E-8:
+ (V(1,2) < 2.230000E0)? 7.942857E-9 * V(1,2) - 1.398257E-8:
+ (V(1,2) < 2.300000E0)? 7.857143E-9 * V(1,2) - 1.379143E-8:
+ (V(1,2) < 2.370000E0)? 7.828571E-9 * V(1,2) - 1.372571E-8:
+ (V(1,2) < 2.440000E0)? 7.671429E-9 * V(1,2) - 1.335329E-8:
+ (V(1,2) < 2.510000E0)? 7.671429E-9 * V(1,2) - 1.335329E-8:
+ (V(1,2) < 2.580000E0)? 7.671429E-9 * V(1,2) - 1.335329E-8:
+ (V(1,2) < 2.650000E0)? 8.000000E-9 * V(1,2) - 1.420100E-8:
+ (V(1,2) < 2.720000E0)? 9.028571E-9 * V(1,2) - 1.692671E-8:
+ (V(1,2) < 2.790000E0)? 9.042857E-9 * V(1,2) - 1.696557E-8:
+ (V(1,2) < 2.860000E0)? 9.042857E-9 * V(1,2) - 1.696557E-8:
+ (V(1,2) < 2.930000E0)? 9.042857E-9 * V(1,2) - 1.696557E-8:
+ (V(1,2) < 3.000000E0)? 1.457143E-8 * V(1,2) - 3.316429E-8:
+ (V(1,2) < 3.070000E0)? 3.200000E-8 * V(1,2) - 8.545000E-8:
+ (V(1,2) < 3.140000E0)? 3.200000E-8 * V(1,2) - 8.545000E-8:
+ (V(1,2) < 3.210000E0)? 3.200000E-8 * V(1,2) - 8.545000E-8:
+ (V(1,2) < 3.280000E0)? 3.200000E-8 * V(1,2) - 8.545000E-8:
+ 1.951000E-8 
.ENDS

************************************* END **************************************


.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-0.5

.SUBCKT NOTUSED N1 N2 N3 N4
* NOTHING HERE: OPEN BETWEEN ALL TERMINALS
.ENDS

