** Circuit for extracting I(OUT)

Rfix DIE OUT 50
Vfix OUT 0 3.3
CComp DIE 0 5.23e-12
VDie DIE 0 PWL(
+ 0 3.3
+ 5.051e-11 3.3
+ 1e-10 3.3
+ 1.5e-10 3.3
+ 2e-10 3.3
+ 2.5e-10 3.3
+ 3e-10 3.3
+ 3.5e-10 3.3
+ 4e-10 3.292
+ 4.5e-10 3.199
+ 5.1e-10 3.128
+ 5.6e-10 3.071
+ 6.1e-10 3.023
+ 6.6e-10 2.982
+ 7.1e-10 2.946
+ 7.6e-10 2.916
+ 8.1e-10 2.889
+ 8.6e-10 2.866
+ 9.1e-10 2.846
+ 9.6e-10 2.828
+ 1.01e-09 2.813
+ 1.06e-09 2.799
+ 1.11e-09 2.787
+ 1.16e-09 2.777
+ 1.21e-09 2.768
+ 1.26e-09 2.76
+ 1.31e-09 2.753
+ 1.36e-09 2.747
+ 1.41e-09 2.741
+ 1.46e-09 2.737
+ 1.52e-09 2.733
+ 1.57e-09 2.729
+ 1.62e-09 2.724
+ 1.67e-09 2.721
+ 1.72e-09 2.72
+ 1.77e-09 2.718
+ 1.82e-09 2.716
+ 1.87e-09 2.714
+ 1.92e-09 2.712
+ 1.97e-09 2.71
+ 2.02e-09 2.708
+ 2.07e-09 2.706
+ 2.12e-09 2.705
+ 2.17e-09 2.704
+ 2.22e-09 2.703
+ 2.27e-09 2.703
+ 2.32e-09 2.702
+ 2.37e-09 2.701
+ 2.42e-09 2.701
+ 2.47e-09 2.7
+ 2.53e-09 2.7
+ 2.58e-09 2.699
+ 2.63e-09 2.699
+ 2.68e-09 2.699
+ 2.73e-09 2.699
+ 2.78e-09 2.699
+ 2.83e-09 2.699
+ 2.88e-09 2.698
+ 2.93e-09 2.698
+ 2.98e-09 2.698
+ 3.03e-09 2.698
+ 3.08e-09 2.698
+ 3.13e-09 2.698
+ 3.18e-09 2.698
+ 3.23e-09 2.698
+ 3.28e-09 2.698
+ 3.33e-09 2.698
+ 3.38e-09 2.698
+ 3.43e-09 2.697
+ 3.48e-09 2.697
+ 3.54e-09 2.697
+ 3.59e-09 2.697
+ 3.64e-09 2.697
+ 3.69e-09 2.697
+ 3.74e-09 2.697
)

.tran 0 3.74e-09
.print tran I(Vdie)
.options NOECHO
.end