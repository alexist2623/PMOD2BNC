********************************************************************************
*
* LTSPICE MODEL FOR IBIS MODEL(S)
* MODELING DATE: 20230619013430
* GENERAETD BY BPRO: http://www.spisim.com
*
* NOTE: ramp data in .ibs model is used in this converted spice model.
*       VT waveform based conversion will yield more accurate result.
*
********************************************************************************


******************************** BEGIN *****************************************
* ORIG. MDL: C:\Jeonghyun\GIT\PMOD2BNC\IBIS\spartan7_v1.3\spartan7\spartan7.ibs;LVCMOS33_S_12_HR;TYP
* TERMINALS: INPUT OUTPUT VCC VSS ENABLE

.SUBCKT LVCMOS33_S_12_HR_TYP NINP NOUT NVCC NVSS NENB

* POWER-ON SOURCE



* INPUT CONTROL
B1 N820 0 V= ((V(NINP) > 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0
B2 N830 0 V= ((V(NINP) < 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0

* RAMP RATE CONTROL
* RISERMP = 1.053709E5 = 1.3722/1.4459n
* FALLRMP = 5.662057E4 = 1.4825/0.8394n

B3 NVCC N850 I= (V(N830) > 0.5)? 0 : V(NVCC, N850) / 5.662057E4
B4 N840 NVSS I= (V(N820) > 0.5)? 0 : V(N840, NVSS) / 1.053709E5
C1 NVCC N850 1F
C2 N840 NVSS 1F
S1 N220 N850 0 N820 SMOD
S2 N840 N220 0 N830 SMOD

G1 N008 NVSS N002 N008 1
G2 NVCC N008 N008 N003 1
R1 N006 NVSS 1
R2 NVCC N006 1

* PU/PD/PC/GC BRANCH
XASRC_PD N002 NVSS N008 N840 LVCMOS33_S_12_HR_PULLDOWN_TYP
XASRC_PU N003 NVCC N850 N008 LVCMOS33_S_12_HR_PULLUP_TYP
XASRC_PC N006 NVCC NVCC N006 LVCMOS33_S_12_HR_POWER_CLAMP_TYP
XASRC_GC N006 NVSS N006 NVSS LVCMOS33_S_12_HR_GND_CLAMP_TYP

* PACKAGE PARASITICS:
ROPKG N001 NOUT 3.345000E-1
COPKG NOUT NVSS 7.200000E-13
LOPKG N005 N001 4.350000E-9
CCOMP N005 NVSS 5.230000E-12

* Voltage Sources for measuring currents
V5 N006 N005 0
V6 N008 N006 0
V7 N220 N008 0
.ENDS

* PU BRANCH
.SUBCKT LVCMOS33_S_12_HR_PULLUP_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -3.300000E0)? 3.786000E-2:
+ (V(1,2) < -3.200000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -3.100000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -3.000000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.900000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.800000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.700000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.600000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.500000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.400000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.300000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.200000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.100000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -2.000000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.900000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.800000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.700000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.600000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.500000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -8.000000E-1)? -0.000000E0 * V(1,2) + 3.786000E-2:
+ (V(1,2) < -7.000000E-1)? -1.910000E-2 * V(1,2) + 2.258000E-2:
+ (V(1,2) < -6.000000E-1)? -7.500000E-3 * V(1,2) + 3.070000E-2:
+ (V(1,2) < -5.000000E-1)? -3.729000E-2 * V(1,2) + 1.282600E-2:
+ (V(1,2) < -4.000000E-1)? -6.070000E-2 * V(1,2) + 1.121000E-3:
+ (V(1,2) < -3.000000E-1)? -4.869200E-2 * V(1,2) + 5.924200E-3:
+ (V(1,2) < -2.000000E-1)? -6.548400E-2 * V(1,2) + 8.866000E-4:
+ (V(1,2) < -1.000000E-1)? -7.053500E-2 * V(1,2) - 1.236000E-4:
+ (V(1,2) < 0.000000E0)? -6.929851E-2 * V(1,2) + 4.936000E-8:
+ (V(1,2) < 1.000000E-1)? -6.506049E-2 * V(1,2) + 4.936000E-8:
+ (V(1,2) < 2.000000E-1)? -6.334000E-2 * V(1,2) - 1.720000E-4:
+ (V(1,2) < 3.000000E-1)? -5.760000E-2 * V(1,2) - 1.320000E-3:
+ (V(1,2) < 4.000000E-1)? -5.300000E-2 * V(1,2) - 2.700000E-3:
+ (V(1,2) < 5.000000E-1)? -4.800000E-2 * V(1,2) - 4.700000E-3:
+ (V(1,2) < 6.000000E-1)? -4.160000E-2 * V(1,2) - 7.900000E-3:
+ (V(1,2) < 7.000000E-1)? -3.990000E-2 * V(1,2) - 8.920000E-3:
+ (V(1,2) < 8.000000E-1)? -3.460000E-2 * V(1,2) - 1.263000E-2:
+ (V(1,2) < 9.000000E-1)? -2.960000E-2 * V(1,2) - 1.663000E-2:
+ (V(1,2) < 1.000000E0)? -2.320000E-2 * V(1,2) - 2.239000E-2:
+ (V(1,2) < 1.100000E0)? -1.920000E-2 * V(1,2) - 2.639000E-2:
+ (V(1,2) < 1.200000E0)? -1.350000E-2 * V(1,2) - 3.266000E-2:
+ (V(1,2) < 1.300000E0)? -9.100000E-3 * V(1,2) - 3.794000E-2:
+ (V(1,2) < 1.400000E0)? -6.000000E-3 * V(1,2) - 4.197000E-2:
+ (V(1,2) < 1.500000E0)? -4.400000E-3 * V(1,2) - 4.421000E-2:
+ (V(1,2) < 1.600000E0)? -3.400000E-3 * V(1,2) - 4.571000E-2:
+ (V(1,2) < 1.700000E0)? -2.900000E-3 * V(1,2) - 4.651000E-2:
+ (V(1,2) < 1.800000E0)? -2.600000E-3 * V(1,2) - 4.702000E-2:
+ (V(1,2) < 1.900000E0)? -2.300000E-3 * V(1,2) - 4.756000E-2:
+ (V(1,2) < 2.000000E0)? -2.100000E-3 * V(1,2) - 4.794000E-2:
+ (V(1,2) < 2.100000E0)? -2.100000E-3 * V(1,2) - 4.794000E-2:
+ (V(1,2) < 2.200000E0)? -1.900000E-3 * V(1,2) - 4.836000E-2:
+ (V(1,2) < 2.300000E0)? -1.800000E-3 * V(1,2) - 4.858000E-2:
+ (V(1,2) < 2.400000E0)? -1.700000E-3 * V(1,2) - 4.881000E-2:
+ (V(1,2) < 2.500000E0)? -9.230000E-2 * V(1,2) + 1.686300E-1:
+ (V(1,2) < 2.600000E0)? -1.300000E-3 * V(1,2) - 5.887000E-2:
+ (V(1,2) < 2.700000E0)? -1.300000E-3 * V(1,2) - 5.887000E-2:
+ (V(1,2) < 2.800000E0)? -1.200000E-3 * V(1,2) - 5.914000E-2:
+ (V(1,2) < 2.900000E0)? -1.200000E-3 * V(1,2) - 5.914000E-2:
+ (V(1,2) < 3.000000E0)? -1.200000E-3 * V(1,2) - 5.914000E-2:
+ (V(1,2) < 3.100000E0)? -1.100000E-3 * V(1,2) - 5.944000E-2:
+ (V(1,2) < 3.200000E0)? -1.100000E-3 * V(1,2) - 5.944000E-2:
+ (V(1,2) < 3.300000E0)? -1.100000E-3 * V(1,2) - 5.944000E-2:
+ (V(1,2) < 3.400000E0)? -1.099000E-3 * V(1,2) - 5.944330E-2:
+ (V(1,2) < 3.500000E0)? -1.187000E-3 * V(1,2) - 5.914410E-2:
+ (V(1,2) < 3.600000E0)? -5.210000E-4 * V(1,2) - 6.147510E-2:
+ (V(1,2) < 3.700000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 3.800000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 3.900000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.000000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.100000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.200000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.300000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.400000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.500000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.600000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.700000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.800000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 4.900000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.000000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.100000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.200000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.300000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.400000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.500000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.600000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.700000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.800000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 5.900000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 6.000000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 6.100000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 6.200000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 6.300000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 6.400000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 6.500000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ (V(1,2) < 6.600000E0)? -0.000000E0 * V(1,2) - 6.335070E-2:
+ -6.335070E-2 
.ENDS

* PD BRANCH
.SUBCKT LVCMOS33_S_12_HR_PULLDOWN_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -3.300000E0)? -4.225000E-2:
+ (V(1,2) < -3.200000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -3.100000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -3.000000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.900000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.800000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.700000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.600000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.500000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.400000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.300000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.200000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.100000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -2.000000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.900000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.800000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.700000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.600000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.500000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -8.000000E-1)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -7.000000E-1)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -6.000000E-1)? -0.000000E0 * V(1,2) - 4.225000E-2:
+ (V(1,2) < -5.000000E-1)? 4.640000E-3 * V(1,2) - 3.946600E-2:
+ (V(1,2) < -4.000000E-1)? 3.610200E-2 * V(1,2) - 2.373500E-2:
+ (V(1,2) < -3.000000E-1)? 9.374500E-2 * V(1,2) - 6.778000E-4:
+ (V(1,2) < -2.000000E-1)? 1.005250E-1 * V(1,2) + 1.356200E-3:
+ (V(1,2) < -1.000000E-1)? 9.777900E-2 * V(1,2) + 8.070000E-4:
+ (V(1,2) < 0.000000E0)? 9.781800E-2 * V(1,2) + 8.109000E-4:
+ (V(1,2) < 1.000000E-1)? 9.111100E-2 * V(1,2) + 8.109000E-4:
+ (V(1,2) < 2.000000E-1)? 6.938000E-2 * V(1,2) + 2.984000E-3:
+ (V(1,2) < 3.000000E-1)? 6.940000E-2 * V(1,2) + 2.980000E-3:
+ (V(1,2) < 4.000000E-1)? 6.940000E-2 * V(1,2) + 2.980000E-3:
+ (V(1,2) < 5.000000E-1)? 6.930000E-2 * V(1,2) + 3.020000E-3:
+ (V(1,2) < 6.000000E-1)? 4.130000E-2 * V(1,2) + 1.702000E-2:
+ (V(1,2) < 7.000000E-1)? 3.380000E-2 * V(1,2) + 2.152000E-2:
+ (V(1,2) < 8.000000E-1)? 3.380000E-2 * V(1,2) + 2.152000E-2:
+ (V(1,2) < 9.000000E-1)? 3.130000E-2 * V(1,2) + 2.352000E-2:
+ (V(1,2) < 1.000000E0)? 6.700000E-3 * V(1,2) + 4.566000E-2:
+ (V(1,2) < 1.100000E0)? 6.700000E-3 * V(1,2) + 4.566000E-2:
+ (V(1,2) < 1.200000E0)? 6.700000E-3 * V(1,2) + 4.566000E-2:
+ (V(1,2) < 1.300000E0)? 5.800000E-3 * V(1,2) + 4.674000E-2:
+ (V(1,2) < 1.400000E0)? 2.700000E-3 * V(1,2) + 5.077000E-2:
+ (V(1,2) < 1.500000E0)? 2.800000E-3 * V(1,2) + 5.063000E-2:
+ (V(1,2) < 1.600000E0)? 2.700000E-3 * V(1,2) + 5.078000E-2:
+ (V(1,2) < 1.700000E0)? 2.000000E-4 * V(1,2) + 5.478000E-2:
+ (V(1,2) < 1.800000E0)? 1.000000E-3 * V(1,2) + 5.342000E-2:
+ (V(1,2) < 1.900000E0)? 1.000000E-3 * V(1,2) + 5.342000E-2:
+ (V(1,2) < 2.000000E0)? 2.400000E-3 * V(1,2) + 5.076000E-2:
+ (V(1,2) < 2.100000E0)? 6.000000E-4 * V(1,2) + 5.436000E-2:
+ (V(1,2) < 2.200000E0)? 1.800000E-3 * V(1,2) + 5.184000E-2:
+ (V(1,2) < 2.300000E0)? -0.000000E0 * V(1,2) + 5.580000E-2:
+ (V(1,2) < 2.400000E0)? 1.200000E-3 * V(1,2) + 5.304000E-2:
+ (V(1,2) < 2.500000E0)? 4.410000E-2 * V(1,2) - 4.992000E-2:
+ (V(1,2) < 2.600000E0)? 3.100000E-3 * V(1,2) + 5.258000E-2:
+ (V(1,2) < 2.700000E0)? 1.100000E-3 * V(1,2) + 5.778000E-2:
+ (V(1,2) < 2.800000E0)? 1.000000E-4 * V(1,2) + 6.048000E-2:
+ (V(1,2) < 2.900000E0)? 6.000000E-4 * V(1,2) + 5.908000E-2:
+ (V(1,2) < 3.000000E0)? 1.000000E-4 * V(1,2) + 6.053000E-2:
+ (V(1,2) < 3.100000E0)? 6.990000E-4 * V(1,2) + 5.873300E-2:
+ (V(1,2) < 3.200000E0)? 2.587000E-3 * V(1,2) + 5.288020E-2:
+ (V(1,2) < 3.300000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 3.400000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 3.500000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 3.600000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 3.700000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 3.800000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 3.900000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.000000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.100000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.200000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.300000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.400000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.500000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.600000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.700000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.800000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 4.900000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.000000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.100000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.200000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.300000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.400000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.500000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.600000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.700000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.800000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 5.900000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 6.000000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 6.100000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 6.200000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 6.300000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 6.400000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 6.500000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ (V(1,2) < 6.600000E0)? -0.000000E0 * V(1,2) + 6.115860E-2:
+ 6.115860E-2 
.ENDS

* PC BRANCH
.SUBCKT LVCMOS33_S_12_HR_POWER_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -3.280000E0)? 3.564000E0:
+ (V(1,2) < -3.240000E0)? -1.550000E0 * V(1,2) - 1.520000E0:
+ (V(1,2) < -3.200000E0)? -1.525000E0 * V(1,2) - 1.439000E0:
+ (V(1,2) < -3.160000E0)? -1.550000E0 * V(1,2) - 1.519000E0:
+ (V(1,2) < -3.120000E0)? -1.525000E0 * V(1,2) - 1.440000E0:
+ (V(1,2) < -3.080000E0)? -1.550000E0 * V(1,2) - 1.518000E0:
+ (V(1,2) < -3.040000E0)? -1.525000E0 * V(1,2) - 1.441000E0:
+ (V(1,2) < -3.000000E0)? -1.550000E0 * V(1,2) - 1.517000E0:
+ (V(1,2) < -2.960000E0)? -1.525000E0 * V(1,2) - 1.442000E0:
+ (V(1,2) < -2.920000E0)? -1.550000E0 * V(1,2) - 1.516000E0:
+ (V(1,2) < -2.880000E0)? -1.525000E0 * V(1,2) - 1.443000E0:
+ (V(1,2) < -2.840000E0)? -1.550000E0 * V(1,2) - 1.515000E0:
+ (V(1,2) < -2.800000E0)? -1.525000E0 * V(1,2) - 1.444000E0:
+ (V(1,2) < -2.760000E0)? -1.525000E0 * V(1,2) - 1.444000E0:
+ (V(1,2) < -2.720000E0)? -1.550000E0 * V(1,2) - 1.513000E0:
+ (V(1,2) < -2.680000E0)? -1.525000E0 * V(1,2) - 1.445000E0:
+ (V(1,2) < -2.640000E0)? -1.550000E0 * V(1,2) - 1.512000E0:
+ (V(1,2) < -2.600000E0)? -1.525000E0 * V(1,2) - 1.446000E0:
+ (V(1,2) < -2.560000E0)? -1.550000E0 * V(1,2) - 1.511000E0:
+ (V(1,2) < -2.520000E0)? -1.525000E0 * V(1,2) - 1.447000E0:
+ (V(1,2) < -2.480000E0)? -1.550000E0 * V(1,2) - 1.510000E0:
+ (V(1,2) < -2.440000E0)? -1.525000E0 * V(1,2) - 1.448000E0:
+ (V(1,2) < -2.400000E0)? -1.550000E0 * V(1,2) - 1.509000E0:
+ (V(1,2) < -2.360000E0)? -1.525000E0 * V(1,2) - 1.449000E0:
+ (V(1,2) < -2.320000E0)? -1.550000E0 * V(1,2) - 1.508000E0:
+ (V(1,2) < -2.280000E0)? -1.525000E0 * V(1,2) - 1.450000E0:
+ (V(1,2) < -2.240000E0)? -1.525000E0 * V(1,2) - 1.450000E0:
+ (V(1,2) < -2.200000E0)? -1.550000E0 * V(1,2) - 1.506000E0:
+ (V(1,2) < -2.160000E0)? -1.525000E0 * V(1,2) - 1.451000E0:
+ (V(1,2) < -2.120000E0)? -1.550000E0 * V(1,2) - 1.505000E0:
+ (V(1,2) < -2.080000E0)? -1.525000E0 * V(1,2) - 1.452000E0:
+ (V(1,2) < -2.040000E0)? -1.550000E0 * V(1,2) - 1.504000E0:
+ (V(1,2) < -2.000000E0)? -1.525000E0 * V(1,2) - 1.453000E0:
+ (V(1,2) < -1.960000E0)? -1.550000E0 * V(1,2) - 1.503000E0:
+ (V(1,2) < -1.920000E0)? -1.525000E0 * V(1,2) - 1.454000E0:
+ (V(1,2) < -1.880000E0)? -1.550000E0 * V(1,2) - 1.502000E0:
+ (V(1,2) < -1.840000E0)? -1.525000E0 * V(1,2) - 1.455000E0:
+ (V(1,2) < -1.800000E0)? -1.525000E0 * V(1,2) - 1.455000E0:
+ (V(1,2) < -1.760000E0)? -1.550000E0 * V(1,2) - 1.500000E0:
+ (V(1,2) < -1.720000E0)? -1.525000E0 * V(1,2) - 1.456000E0:
+ (V(1,2) < -1.680000E0)? -1.550000E0 * V(1,2) - 1.499000E0:
+ (V(1,2) < -1.640000E0)? -1.525000E0 * V(1,2) - 1.457000E0:
+ (V(1,2) < -1.600000E0)? -1.532500E0 * V(1,2) - 1.469300E0:
+ (V(1,2) < -1.560000E0)? -1.535000E0 * V(1,2) - 1.473300E0:
+ (V(1,2) < -1.520000E0)? -1.532500E0 * V(1,2) - 1.469400E0:
+ (V(1,2) < -1.480000E0)? -1.532500E0 * V(1,2) - 1.469400E0:
+ (V(1,2) < -1.440000E0)? -1.530000E0 * V(1,2) - 1.465700E0:
+ (V(1,2) < -1.400000E0)? -1.532500E0 * V(1,2) - 1.469300E0:
+ (V(1,2) < -1.360000E0)? -1.530000E0 * V(1,2) - 1.465800E0:
+ (V(1,2) < -1.320000E0)? -1.492500E0 * V(1,2) - 1.414800E0:
+ (V(1,2) < -1.280000E0)? -1.465000E0 * V(1,2) - 1.378500E0:
+ (V(1,2) < -1.240000E0)? -1.465000E0 * V(1,2) - 1.378500E0:
+ (V(1,2) < -1.200000E0)? -1.462500E0 * V(1,2) - 1.375400E0:
+ (V(1,2) < -1.160000E0)? -1.465000E0 * V(1,2) - 1.378400E0:
+ (V(1,2) < -1.120000E0)? -1.367500E0 * V(1,2) - 1.265300E0:
+ (V(1,2) < -1.080000E0)? -1.290000E0 * V(1,2) - 1.178500E0:
+ (V(1,2) < -1.040000E0)? -1.292500E0 * V(1,2) - 1.181200E0:
+ (V(1,2) < -1.000000E0)? -1.125000E0 * V(1,2) - 1.007000E0:
+ (V(1,2) < -9.600000E-1)? -9.245000E-1 * V(1,2) - 8.065000E-1:
+ (V(1,2) < -9.200000E-1)? -6.370000E-1 * V(1,2) - 5.305000E-1:
+ (V(1,2) < -8.800000E-1)? -3.540000E-1 * V(1,2) - 2.701400E-1:
+ (V(1,2) < -8.400000E-1)? -2.055000E-1 * V(1,2) - 1.394600E-1:
+ (V(1,2) < -8.000000E-1)? -1.277500E-1 * V(1,2) - 7.415000E-2:
+ (V(1,2) < -7.600000E-1)? -8.875000E-2 * V(1,2) - 4.295000E-2:
+ (V(1,2) < -7.200000E-1)? -8.425000E-2 * V(1,2) - 3.953000E-2:
+ (V(1,2) < -6.800000E-1)? -8.450000E-2 * V(1,2) - 3.971000E-2:
+ (V(1,2) < -6.400000E-1)? -8.450000E-2 * V(1,2) - 3.971000E-2:
+ (V(1,2) < -6.000000E-1)? -8.450000E-2 * V(1,2) - 3.971000E-2:
+ (V(1,2) < -5.600000E-1)? -5.177500E-2 * V(1,2) - 2.007500E-2:
+ (V(1,2) < -5.200000E-1)? -4.837500E-2 * V(1,2) - 1.817100E-2:
+ (V(1,2) < -4.800000E-1)? -4.835000E-2 * V(1,2) - 1.815800E-2:
+ (V(1,2) < -4.400000E-1)? -4.835000E-2 * V(1,2) - 1.815800E-2:
+ (V(1,2) < -4.000000E-1)? -4.835000E-2 * V(1,2) - 1.815800E-2:
+ (V(1,2) < -3.600000E-1)? -9.712500E-3 * V(1,2) - 2.703000E-3:
+ (V(1,2) < -3.200000E-1)? -5.767500E-3 * V(1,2) - 1.282800E-3:
+ (V(1,2) < -2.800000E-1)? -5.765000E-3 * V(1,2) - 1.282000E-3:
+ (V(1,2) < -2.400000E-1)? -5.767500E-3 * V(1,2) - 1.282700E-3:
+ (V(1,2) < -2.000000E-1)? -2.419775E-3 * V(1,2) - 4.792460E-4:
+ (V(1,2) < -1.600000E-1)? -5.147500E-5 * V(1,2) - 5.586000E-6:
+ (V(1,2) < -1.200000E-1)? -5.149000E-5 * V(1,2) - 5.588400E-6:
+ (V(1,2) < -8.000000E-2)? -1.278325E-5 * V(1,2) - 9.435900E-7:
+ (V(1,2) < -4.000000E-2)? -1.242250E-6 * V(1,2) - 2.031000E-8:
+ (V(1,2) < 0.000000E0)? -2.440000E-7 * V(1,2) + 1.962000E-8:
+ 1.962000E-8 
.ENDS

* GC BRANCH
.SUBCKT LVCMOS33_S_12_HR_GND_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -3.300000E0)? -3.592000E0:
+ (V(1,2) < -3.230000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -3.160000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -3.090000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -3.020000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -2.950000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -2.880000E0)? 1.528571E0 * V(1,2) + 1.452286E0:
+ (V(1,2) < -2.810000E0)? 1.514286E0 * V(1,2) + 1.411143E0:
+ (V(1,2) < -2.740000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.670000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.600000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.530000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.460000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.390000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.320000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.250000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.180000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.110000E0)? 1.528571E0 * V(1,2) + 1.451286E0:
+ (V(1,2) < -2.040000E0)? 1.514286E0 * V(1,2) + 1.421143E0:
+ (V(1,2) < -1.970000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.900000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.830000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.760000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.690000E0)? 1.528571E0 * V(1,2) + 1.450286E0:
+ (V(1,2) < -1.620000E0)? 1.514286E0 * V(1,2) + 1.426143E0:
+ (V(1,2) < -1.550000E0)? 1.498571E0 * V(1,2) + 1.400686E0:
+ (V(1,2) < -1.480000E0)? 1.500000E0 * V(1,2) + 1.402900E0:
+ (V(1,2) < -1.410000E0)? 1.500000E0 * V(1,2) + 1.402900E0:
+ (V(1,2) < -1.340000E0)? 1.501429E0 * V(1,2) + 1.404914E0:
+ (V(1,2) < -1.270000E0)? 1.457143E0 * V(1,2) + 1.345571E0:
+ (V(1,2) < -1.200000E0)? 1.201429E0 * V(1,2) + 1.020814E0:
+ (V(1,2) < -1.130000E0)? 1.200000E0 * V(1,2) + 1.019100E0:
+ (V(1,2) < -1.060000E0)? 1.201429E0 * V(1,2) + 1.020714E0:
+ (V(1,2) < -9.900000E-1)? 1.200000E0 * V(1,2) + 1.019200E0:
+ (V(1,2) < -9.200000E-1)? 1.092857E0 * V(1,2) + 9.131286E-1:
+ (V(1,2) < -8.500000E-1)? 4.321429E-1 * V(1,2) + 3.052714E-1:
+ (V(1,2) < -7.800000E-1)? 2.414286E-1 * V(1,2) + 1.431643E-1:
+ (V(1,2) < -7.100000E-1)? 1.680000E-1 * V(1,2) + 8.589000E-2:
+ (V(1,2) < -6.400000E-1)? 1.680000E-1 * V(1,2) + 8.589000E-2:
+ (V(1,2) < -5.700000E-1)? 1.198571E-1 * V(1,2) + 5.507857E-2:
+ (V(1,2) < -5.000000E-1)? 9.605714E-2 * V(1,2) + 4.151257E-2:
+ (V(1,2) < -4.300000E-1)? 7.432857E-2 * V(1,2) + 3.064829E-2:
+ (V(1,2) < -3.600000E-1)? 1.554429E-2 * V(1,2) + 5.371043E-3:
+ (V(1,2) < -2.900000E-1)? 2.747857E-3 * V(1,2) + 7.643286E-4:
+ (V(1,2) < -2.200000E-1)? 3.692286E-4 * V(1,2) + 7.452629E-5:
+ (V(1,2) < -1.500000E-1)? 9.002714E-5 * V(1,2) + 1.310197E-5:
+ (V(1,2) < -8.000000E-2)? 5.286714E-6 * V(1,2) + 3.909071E-7:
+ (V(1,2) < -1.000000E-2)? 2.521429E-7 * V(1,2) - 1.185857E-8:
+ (V(1,2) < 6.000000E-2)? 3.014286E-8 * V(1,2) - 1.407857E-8:
+ (V(1,2) < 1.300000E-1)? 1.300000E-8 * V(1,2) - 1.305000E-8:
+ (V(1,2) < 2.000000E-1)? 8.714286E-9 * V(1,2) - 1.249286E-8:
+ (V(1,2) < 2.700000E-1)? 6.857143E-9 * V(1,2) - 1.212143E-8:
+ (V(1,2) < 3.400000E-1)? 6.342857E-9 * V(1,2) - 1.198257E-8:
+ (V(1,2) < 4.100000E-1)? 5.885714E-9 * V(1,2) - 1.182714E-8:
+ (V(1,2) < 4.800000E-1)? 5.842857E-9 * V(1,2) - 1.180957E-8:
+ (V(1,2) < 5.500000E-1)? 5.600000E-9 * V(1,2) - 1.169300E-8:
+ (V(1,2) < 6.200000E-1)? 5.542857E-9 * V(1,2) - 1.166157E-8:
+ (V(1,2) < 6.900000E-1)? 5.428571E-9 * V(1,2) - 1.159071E-8:
+ (V(1,2) < 7.600000E-1)? 5.414286E-9 * V(1,2) - 1.158086E-8:
+ (V(1,2) < 8.300000E-1)? 5.400000E-9 * V(1,2) - 1.157000E-8:
+ (V(1,2) < 9.000000E-1)? 5.385714E-9 * V(1,2) - 1.155814E-8:
+ (V(1,2) < 9.700000E-1)? 5.371429E-9 * V(1,2) - 1.154529E-8:
+ (V(1,2) < 1.040000E0)? 5.428571E-9 * V(1,2) - 1.160071E-8:
+ (V(1,2) < 1.110000E0)? 5.371429E-9 * V(1,2) - 1.154129E-8:
+ (V(1,2) < 1.180000E0)? 5.442857E-9 * V(1,2) - 1.162057E-8:
+ (V(1,2) < 1.250000E0)? 5.214286E-9 * V(1,2) - 1.135086E-8:
+ (V(1,2) < 1.320000E0)? 5.014286E-9 * V(1,2) - 1.110086E-8:
+ (V(1,2) < 1.390000E0)? 5.128571E-9 * V(1,2) - 1.125171E-8:
+ (V(1,2) < 1.460000E0)? 5.500000E-9 * V(1,2) - 1.176800E-8:
+ (V(1,2) < 1.530000E0)? 7.700000E-9 * V(1,2) - 1.498000E-8:
+ (V(1,2) < 1.600000E0)? 9.685714E-9 * V(1,2) - 1.801814E-8:
+ (V(1,2) < 1.670000E0)? 1.100000E-8 * V(1,2) - 2.012100E-8:
+ (V(1,2) < 1.740000E0)? 1.142857E-8 * V(1,2) - 2.083671E-8:
+ (V(1,2) < 1.810000E0)? 9.262857E-9 * V(1,2) - 1.706837E-8:
+ (V(1,2) < 1.880000E0)? 1.195571E-8 * V(1,2) - 2.194244E-8:
+ (V(1,2) < 1.950000E0)? 1.421000E-8 * V(1,2) - 2.618050E-8:
+ (V(1,2) < 2.020000E0)? 7.828571E-9 * V(1,2) - 1.373671E-8:
+ (V(1,2) < 2.090000E0)? 7.071429E-9 * V(1,2) - 1.220729E-8:
+ (V(1,2) < 2.160000E0)? 8.685714E-9 * V(1,2) - 1.558114E-8:
+ (V(1,2) < 2.230000E0)? 8.057143E-9 * V(1,2) - 1.422343E-8:
+ (V(1,2) < 2.300000E0)? 7.571429E-9 * V(1,2) - 1.314029E-8:
+ (V(1,2) < 2.370000E0)? 7.614286E-9 * V(1,2) - 1.323886E-8:
+ (V(1,2) < 2.440000E0)? 7.814286E-9 * V(1,2) - 1.371286E-8:
+ (V(1,2) < 2.510000E0)? 7.828571E-9 * V(1,2) - 1.374771E-8:
+ (V(1,2) < 2.580000E0)? 7.828571E-9 * V(1,2) - 1.374771E-8:
+ (V(1,2) < 2.650000E0)? 8.128571E-9 * V(1,2) - 1.452171E-8:
+ (V(1,2) < 2.720000E0)? 8.885714E-9 * V(1,2) - 1.652814E-8:
+ (V(1,2) < 2.790000E0)? 8.900000E-9 * V(1,2) - 1.656700E-8:
+ (V(1,2) < 2.860000E0)? 8.885714E-9 * V(1,2) - 1.652714E-8:
+ (V(1,2) < 2.930000E0)? 8.900000E-9 * V(1,2) - 1.656800E-8:
+ (V(1,2) < 3.000000E0)? 1.044286E-8 * V(1,2) - 2.108857E-8:
+ (V(1,2) < 3.070000E0)? 1.771429E-8 * V(1,2) - 4.290286E-8:
+ (V(1,2) < 3.140000E0)? 3.757143E-8 * V(1,2) - 1.038643E-7:
+ (V(1,2) < 3.210000E0)? 3.771429E-8 * V(1,2) - 1.043129E-7:
+ (V(1,2) < 3.280000E0)? 3.771429E-8 * V(1,2) - 1.043129E-7:
+ 1.939000E-8 
.ENDS

************************************* END **************************************


.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-0.5

.SUBCKT NOTUSED N1 N2 N3 N4
* NOTHING HERE: OPEN BETWEEN ALL TERMINALS
.ENDS

