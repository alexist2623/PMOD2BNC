

.subckt TL_SL1 1 2 ngnd length=0.150081


WTL1 1 ngnd 2 ngnd n=1 RLGCfile=G6Q2.rlc l='length'



.ends TL_SL1
