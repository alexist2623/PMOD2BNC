

.subckt resistorPack_850 G1 S1 S2 S3 S4 S5 S6 S7


R1 S1 G1 50
R2 S2 G1 50
R3 S3 G1 50
R4 S4 G1 50
R5 S5 G1 50
R6 S6 G1 50
R7 S7 G1 50


.ends resistorPack_850
