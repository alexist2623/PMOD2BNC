********************************************************************************
*
* LTSPICE MODEL FOR IBIS MODEL(S)
* MODELING DATE: 20230603112723
* GENERAETD BY BPRO: http://www.spisim.com
*
* NOTE: ramp data in .ibs model is used in this converted spice model.
*       VT waveform based conversion will yield more accurate result.
*
********************************************************************************


******************************** BEGIN *****************************************
* ORIG. MDL: C:\Jeonghyun\GIT\PMOD2BNC\IBIS\spartan7_v1.3\spartan7\spartan7.ibs;HSTL_II_F_HR_IN50;TYP
* TERMINALS: INPUT OUTPUT VCC VSS ENABLE

.SUBCKT HSTL_II_F_HR_IN50_TYP NINP NOUT NVCC NVSS NENB

* POWER-ON SOURCE



* INPUT CONTROL
B1 N820 0 V= ((V(NINP) > 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0
B2 N830 0 V= ((V(NINP) < 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0

* RAMP RATE CONTROL
* RISERMP = 3.005958E4 = 0.5539/0.1665n
* FALLRMP = 3.456172E4 = 0.5590/0.1932n

B3 NVCC N850 I= (V(N830) > 0.5)? 0 : V(NVCC, N850) / 3.456172E4
B4 N840 NVSS I= (V(N820) > 0.5)? 0 : V(N840, NVSS) / 3.005958E4
C1 NVCC N850 1F
C2 N840 NVSS 1F
S1 N220 N850 0 N820 SMOD
S2 N840 N220 0 N830 SMOD

G1 N008 NVSS N002 N008 1
G2 NVCC N008 N008 N003 1
R1 N006 NVSS 1
R2 NVCC N006 1

* PU/PD/PC/GC BRANCH
XASRC_PD N002 NVSS N008 N840 HSTL_II_F_HR_IN50_PULLDOWN_TYP
XASRC_PU N003 NVCC N850 N008 HSTL_II_F_HR_IN50_PULLUP_TYP
XASRC_PC N006 NVCC NVCC N006 HSTL_II_F_HR_IN50_POWER_CLAMP_TYP
XASRC_GC N006 NVSS N006 NVSS HSTL_II_F_HR_IN50_GND_CLAMP_TYP

* PACKAGE PARASITICS:
ROPKG N001 NOUT 3.345000E-1
COPKG NOUT NVSS 7.200000E-13
LOPKG N005 N001 4.350000E-9
CCOMP N005 NVSS 7.690000E-12

* Voltage Sources for measuring currents
V5 N006 N005 0
V6 N008 N006 0
V7 N220 N008 0
.ENDS

* PU BRANCH
.SUBCKT HSTL_II_F_HR_IN50_PULLUP_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -1.500000E0)? 6.717000E-2:
+ (V(1,2) < -1.450000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.350000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.250000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.150000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.050000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -9.500000E-1)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -8.500000E-1)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -8.000000E-1)? -0.000000E0 * V(1,2) + 6.717000E-2:
+ (V(1,2) < -7.500000E-1)? -2.986000E-2 * V(1,2) + 4.328200E-2:
+ (V(1,2) < -7.000000E-1)? -4.876000E-2 * V(1,2) + 2.910700E-2:
+ (V(1,2) < -6.500000E-1)? -6.624000E-2 * V(1,2) + 1.687100E-2:
+ (V(1,2) < -6.000000E-1)? -8.302600E-2 * V(1,2) + 5.960100E-3:
+ (V(1,2) < -5.500000E-1)? -9.417200E-2 * V(1,2) - 7.275000E-4:
+ (V(1,2) < -5.000000E-1)? -9.794400E-2 * V(1,2) - 2.802100E-3:
+ (V(1,2) < -4.500000E-1)? -9.794000E-2 * V(1,2) - 2.800100E-3:
+ (V(1,2) < -4.000000E-1)? -9.712400E-2 * V(1,2) - 2.432900E-3:
+ (V(1,2) < -3.500000E-1)? -9.584200E-2 * V(1,2) - 1.920100E-3:
+ (V(1,2) < -3.000000E-1)? -9.451800E-2 * V(1,2) - 1.456700E-3:
+ (V(1,2) < -2.500000E-1)? -9.338000E-2 * V(1,2) - 1.115300E-3:
+ (V(1,2) < -2.000000E-1)? -9.179600E-2 * V(1,2) - 7.193000E-4:
+ (V(1,2) < -1.500000E-1)? -9.039800E-2 * V(1,2) - 4.397000E-4:
+ (V(1,2) < -1.000000E-1)? -8.908000E-2 * V(1,2) - 2.420000E-4:
+ (V(1,2) < -5.000000E-2)? -8.746000E-2 * V(1,2) - 8.000000E-5:
+ (V(1,2) < 0.000000E0)? -8.586001E-2 * V(1,2) - 3.960000E-10:
+ (V(1,2) < 5.000000E-2)? -8.331999E-2 * V(1,2) - 3.960000E-10:
+ (V(1,2) < 1.000000E-1)? -7.988000E-2 * V(1,2) - 1.720000E-4:
+ (V(1,2) < 1.500000E-1)? -7.640000E-2 * V(1,2) - 5.200000E-4:
+ (V(1,2) < 2.000000E-1)? -7.280000E-2 * V(1,2) - 1.060000E-3:
+ (V(1,2) < 2.500000E-1)? -6.920000E-2 * V(1,2) - 1.780000E-3:
+ (V(1,2) < 3.000000E-1)? -6.540000E-2 * V(1,2) - 2.730000E-3:
+ (V(1,2) < 3.500000E-1)? -6.160000E-2 * V(1,2) - 3.870000E-3:
+ (V(1,2) < 4.000000E-1)? -5.800000E-2 * V(1,2) - 5.130000E-3:
+ (V(1,2) < 4.500000E-1)? -5.380000E-2 * V(1,2) - 6.810000E-3:
+ (V(1,2) < 5.000000E-1)? -5.000000E-2 * V(1,2) - 8.520000E-3:
+ (V(1,2) < 5.500000E-1)? -4.580000E-2 * V(1,2) - 1.062000E-2:
+ (V(1,2) < 6.000000E-1)? -4.180000E-2 * V(1,2) - 1.282000E-2:
+ (V(1,2) < 6.500000E-1)? -3.760000E-2 * V(1,2) - 1.534000E-2:
+ (V(1,2) < 7.000000E-1)? -3.340000E-2 * V(1,2) - 1.807000E-2:
+ (V(1,2) < 7.500000E-1)? -2.940000E-2 * V(1,2) - 2.087000E-2:
+ (V(1,2) < 8.000000E-1)? -2.520000E-2 * V(1,2) - 2.402000E-2:
+ (V(1,2) < 8.500000E-1)? -2.120000E-2 * V(1,2) - 2.722000E-2:
+ (V(1,2) < 9.000000E-1)? -1.760000E-2 * V(1,2) - 3.028000E-2:
+ (V(1,2) < 9.500000E-1)? -1.440000E-2 * V(1,2) - 3.316000E-2:
+ (V(1,2) < 1.000000E0)? -1.180000E-2 * V(1,2) - 3.563000E-2:
+ (V(1,2) < 1.050000E0)? -1.000000E-2 * V(1,2) - 3.743000E-2:
+ (V(1,2) < 1.100000E0)? -8.600000E-3 * V(1,2) - 3.890000E-2:
+ (V(1,2) < 1.150000E0)? -7.600000E-3 * V(1,2) - 4.000000E-2:
+ (V(1,2) < 1.200000E0)? -6.600000E-3 * V(1,2) - 4.115000E-2:
+ (V(1,2) < 1.250000E0)? -6.200000E-3 * V(1,2) - 4.163000E-2:
+ (V(1,2) < 1.300000E0)? -5.600000E-3 * V(1,2) - 4.238000E-2:
+ (V(1,2) < 1.350000E0)? -5.400000E-3 * V(1,2) - 4.264000E-2:
+ (V(1,2) < 1.400000E0)? -5.000000E-3 * V(1,2) - 4.318000E-2:
+ (V(1,2) < 1.450000E0)? -4.600000E-3 * V(1,2) - 4.374000E-2:
+ (V(1,2) < 1.500000E0)? -4.600000E-3 * V(1,2) - 4.374000E-2:
+ (V(1,2) < 1.550000E0)? -4.200000E-3 * V(1,2) - 4.434000E-2:
+ (V(1,2) < 1.600000E0)? -4.200000E-3 * V(1,2) - 4.434000E-2:
+ (V(1,2) < 1.650000E0)? -3.998000E-3 * V(1,2) - 4.466320E-2:
+ (V(1,2) < 1.700000E0)? -3.986000E-3 * V(1,2) - 4.468300E-2:
+ (V(1,2) < 1.750000E0)? -3.722000E-3 * V(1,2) - 4.513180E-2:
+ (V(1,2) < 1.800000E0)? -3.390000E-3 * V(1,2) - 4.571280E-2:
+ (V(1,2) < 1.850000E0)? -2.432000E-3 * V(1,2) - 4.743720E-2:
+ (V(1,2) < 1.900000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 1.950000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.000000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.050000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.100000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.150000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.200000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.250000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.300000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.350000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.400000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.450000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.500000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.550000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.600000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.650000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.700000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.750000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.800000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.850000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.900000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 2.950000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ (V(1,2) < 3.000000E0)? -0.000000E0 * V(1,2) - 5.193640E-2:
+ -5.193640E-2 
.ENDS

* PD BRANCH
.SUBCKT HSTL_II_F_HR_IN50_PULLDOWN_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -1.500000E0)? -4.122000E-2:
+ (V(1,2) < -1.450000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.350000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.250000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.150000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.050000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -9.500000E-1)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -8.500000E-1)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -8.000000E-1)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -7.500000E-1)? -0.000000E0 * V(1,2) - 4.122000E-2:
+ (V(1,2) < -7.000000E-1)? 2.000000E-4 * V(1,2) - 4.107000E-2:
+ (V(1,2) < -6.500000E-1)? 2.600000E-3 * V(1,2) - 3.939000E-2:
+ (V(1,2) < -6.000000E-1)? 5.600000E-3 * V(1,2) - 3.744000E-2:
+ (V(1,2) < -5.500000E-1)? 1.254000E-2 * V(1,2) - 3.327600E-2:
+ (V(1,2) < -5.000000E-1)? 2.444000E-2 * V(1,2) - 2.673100E-2:
+ (V(1,2) < -4.500000E-1)? 4.260000E-2 * V(1,2) - 1.765100E-2:
+ (V(1,2) < -4.000000E-1)? 6.128200E-2 * V(1,2) - 9.244100E-3:
+ (V(1,2) < -3.500000E-1)? 7.381000E-2 * V(1,2) - 4.232900E-3:
+ (V(1,2) < -3.000000E-1)? 7.923200E-2 * V(1,2) - 2.335200E-3:
+ (V(1,2) < -2.500000E-1)? 8.199000E-2 * V(1,2) - 1.507800E-3:
+ (V(1,2) < -2.000000E-1)? 8.392200E-2 * V(1,2) - 1.024800E-3:
+ (V(1,2) < -1.500000E-1)? 8.598600E-2 * V(1,2) - 6.120000E-4:
+ (V(1,2) < -1.000000E-1)? 8.787800E-2 * V(1,2) - 3.282000E-4:
+ (V(1,2) < -5.000000E-2)? 9.006000E-2 * V(1,2) - 1.100000E-4:
+ (V(1,2) < 0.000000E0)? 9.226000E-2 * V(1,2) + 1.710000E-10:
+ (V(1,2) < 5.000000E-2)? 9.076000E-2 * V(1,2) + 1.710000E-10:
+ (V(1,2) < 1.000000E-1)? 8.560000E-2 * V(1,2) + 2.580000E-4:
+ (V(1,2) < 1.500000E-1)? 8.064000E-2 * V(1,2) + 7.540000E-4:
+ (V(1,2) < 2.000000E-1)? 7.540000E-2 * V(1,2) + 1.540000E-3:
+ (V(1,2) < 2.500000E-1)? 7.080000E-2 * V(1,2) + 2.460000E-3:
+ (V(1,2) < 3.000000E-1)? 6.600000E-2 * V(1,2) + 3.660000E-3:
+ (V(1,2) < 3.500000E-1)? 6.120000E-2 * V(1,2) + 5.100000E-3:
+ (V(1,2) < 4.000000E-1)? 5.680000E-2 * V(1,2) + 6.640000E-3:
+ (V(1,2) < 4.500000E-1)? 5.220000E-2 * V(1,2) + 8.480000E-3:
+ (V(1,2) < 5.000000E-1)? 4.800000E-2 * V(1,2) + 1.037000E-2:
+ (V(1,2) < 5.500000E-1)? 4.360000E-2 * V(1,2) + 1.257000E-2:
+ (V(1,2) < 6.000000E-1)? 3.940000E-2 * V(1,2) + 1.488000E-2:
+ (V(1,2) < 6.500000E-1)? 3.520000E-2 * V(1,2) + 1.740000E-2:
+ (V(1,2) < 7.000000E-1)? 3.120000E-2 * V(1,2) + 2.000000E-2:
+ (V(1,2) < 7.500000E-1)? 2.720000E-2 * V(1,2) + 2.280000E-2:
+ (V(1,2) < 8.000000E-1)? 2.340000E-2 * V(1,2) + 2.565000E-2:
+ (V(1,2) < 8.500000E-1)? 1.980000E-2 * V(1,2) + 2.853000E-2:
+ (V(1,2) < 9.000000E-1)? 1.640000E-2 * V(1,2) + 3.142000E-2:
+ (V(1,2) < 9.500000E-1)? 1.340000E-2 * V(1,2) + 3.412000E-2:
+ (V(1,2) < 1.000000E0)? 1.080000E-2 * V(1,2) + 3.659000E-2:
+ (V(1,2) < 1.050000E0)? 8.400000E-3 * V(1,2) + 3.899000E-2:
+ (V(1,2) < 1.100000E0)? 6.600000E-3 * V(1,2) + 4.088000E-2:
+ (V(1,2) < 1.150000E0)? 5.000000E-3 * V(1,2) + 4.264000E-2:
+ (V(1,2) < 1.200000E0)? 3.600000E-3 * V(1,2) + 4.425000E-2:
+ (V(1,2) < 1.250000E0)? 3.000000E-3 * V(1,2) + 4.497000E-2:
+ (V(1,2) < 1.300000E0)? 2.200000E-3 * V(1,2) + 4.597000E-2:
+ (V(1,2) < 1.350000E0)? 1.800000E-3 * V(1,2) + 4.649000E-2:
+ (V(1,2) < 1.400000E0)? 1.600000E-3 * V(1,2) + 4.676000E-2:
+ (V(1,2) < 1.450000E0)? 1.200000E-3 * V(1,2) + 4.732000E-2:
+ (V(1,2) < 1.500000E0)? 1.200000E-3 * V(1,2) + 4.732000E-2:
+ (V(1,2) < 1.550000E0)? 1.000000E-3 * V(1,2) + 4.762000E-2:
+ (V(1,2) < 1.600000E0)? 1.000000E-3 * V(1,2) + 4.762000E-2:
+ (V(1,2) < 1.650000E0)? 1.000000E-3 * V(1,2) + 4.762000E-2:
+ (V(1,2) < 1.700000E0)? 7.980000E-4 * V(1,2) + 4.795330E-2:
+ (V(1,2) < 1.750000E0)? 7.960000E-4 * V(1,2) + 4.795670E-2:
+ (V(1,2) < 1.800000E0)? 5.800000E-4 * V(1,2) + 4.833470E-2:
+ (V(1,2) < 1.850000E0)? 7.180000E-4 * V(1,2) + 4.808630E-2:
+ (V(1,2) < 1.900000E0)? 8.420000E-4 * V(1,2) + 4.785690E-2:
+ (V(1,2) < 1.950000E0)? 3.240000E-4 * V(1,2) + 4.884110E-2:
+ (V(1,2) < 2.000000E0)? 3.400000E-4 * V(1,2) + 4.880990E-2:
+ (V(1,2) < 2.050000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.100000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.150000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.200000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.250000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.300000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.350000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.400000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.450000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.500000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.550000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.600000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.650000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.700000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.750000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.800000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.850000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.900000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 2.950000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ (V(1,2) < 3.000000E0)? -0.000000E0 * V(1,2) + 4.948990E-2:
+ 4.948990E-2 
.ENDS

* PC BRANCH
.SUBCKT HSTL_II_F_HR_IN50_POWER_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -1.500000E0)? 8.278000E-1:
+ (V(1,2) < -1.480000E0)? -1.535000E0 * V(1,2) - 1.474700E0:
+ (V(1,2) < -1.460000E0)? -1.535000E0 * V(1,2) - 1.474700E0:
+ (V(1,2) < -1.440000E0)? -1.535000E0 * V(1,2) - 1.474700E0:
+ (V(1,2) < -1.420000E0)? -1.540000E0 * V(1,2) - 1.481900E0:
+ (V(1,2) < -1.400000E0)? -1.530000E0 * V(1,2) - 1.467700E0:
+ (V(1,2) < -1.380000E0)? -1.530000E0 * V(1,2) - 1.467700E0:
+ (V(1,2) < -1.360000E0)? -1.525000E0 * V(1,2) - 1.460800E0:
+ (V(1,2) < -1.340000E0)? -1.515000E0 * V(1,2) - 1.447200E0:
+ (V(1,2) < -1.320000E0)? -1.515000E0 * V(1,2) - 1.447200E0:
+ (V(1,2) < -1.300000E0)? -1.505000E0 * V(1,2) - 1.434000E0:
+ (V(1,2) < -1.280000E0)? -1.495000E0 * V(1,2) - 1.421000E0:
+ (V(1,2) < -1.260000E0)? -1.490000E0 * V(1,2) - 1.414600E0:
+ (V(1,2) < -1.240000E0)? -1.480000E0 * V(1,2) - 1.402000E0:
+ (V(1,2) < -1.220000E0)? -1.470000E0 * V(1,2) - 1.389600E0:
+ (V(1,2) < -1.200000E0)? -1.455000E0 * V(1,2) - 1.371300E0:
+ (V(1,2) < -1.180000E0)? -1.445000E0 * V(1,2) - 1.359300E0:
+ (V(1,2) < -1.160000E0)? -1.425000E0 * V(1,2) - 1.335700E0:
+ (V(1,2) < -1.140000E0)? -1.410000E0 * V(1,2) - 1.318300E0:
+ (V(1,2) < -1.120000E0)? -1.385000E0 * V(1,2) - 1.289800E0:
+ (V(1,2) < -1.100000E0)? -1.360000E0 * V(1,2) - 1.261800E0:
+ (V(1,2) < -1.080000E0)? -1.330000E0 * V(1,2) - 1.228800E0:
+ (V(1,2) < -1.060000E0)? -1.290000E0 * V(1,2) - 1.185600E0:
+ (V(1,2) < -1.040000E0)? -1.245000E0 * V(1,2) - 1.137900E0:
+ (V(1,2) < -1.020000E0)? -1.190000E0 * V(1,2) - 1.080700E0:
+ (V(1,2) < -1.000000E0)? -1.115000E0 * V(1,2) - 1.004200E0:
+ (V(1,2) < -9.800000E-1)? -1.027000E0 * V(1,2) - 9.162000E-1:
+ (V(1,2) < -9.600000E-1)? -9.185000E-1 * V(1,2) - 8.098700E-1:
+ (V(1,2) < -9.400000E-1)? -7.890000E-1 * V(1,2) - 6.855500E-1:
+ (V(1,2) < -9.200000E-1)? -6.450000E-1 * V(1,2) - 5.501900E-1:
+ (V(1,2) < -9.000000E-1)? -4.990000E-1 * V(1,2) - 4.158700E-1:
+ (V(1,2) < -8.800000E-1)? -3.690000E-1 * V(1,2) - 2.988700E-1:
+ (V(1,2) < -8.600000E-1)? -2.650000E-1 * V(1,2) - 2.073500E-1:
+ (V(1,2) < -8.400000E-1)? -1.930000E-1 * V(1,2) - 1.454300E-1:
+ (V(1,2) < -8.200000E-1)? -1.460000E-1 * V(1,2) - 1.059500E-1:
+ (V(1,2) < -8.000000E-1)? -1.165000E-1 * V(1,2) - 8.176000E-2:
+ (V(1,2) < -7.800000E-1)? -9.830000E-2 * V(1,2) - 6.720000E-2:
+ (V(1,2) < -7.600000E-1)? -8.530000E-2 * V(1,2) - 5.706000E-2:
+ (V(1,2) < -7.400000E-1)? -7.525000E-2 * V(1,2) - 4.942200E-2:
+ (V(1,2) < -7.200000E-1)? -6.650000E-2 * V(1,2) - 4.294700E-2:
+ (V(1,2) < -7.000000E-1)? -5.810000E-2 * V(1,2) - 3.689900E-2:
+ (V(1,2) < -6.800000E-1)? -4.955000E-2 * V(1,2) - 3.091400E-2:
+ (V(1,2) < -6.600000E-1)? -4.075000E-2 * V(1,2) - 2.493000E-2:
+ (V(1,2) < -6.400000E-1)? -3.195000E-2 * V(1,2) - 1.912200E-2:
+ (V(1,2) < -6.200000E-1)? -2.366500E-2 * V(1,2) - 1.381960E-2:
+ (V(1,2) < -6.000000E-1)? -1.642000E-2 * V(1,2) - 9.327700E-3:
+ (V(1,2) < -5.800000E-1)? -1.072500E-2 * V(1,2) - 5.910700E-3:
+ (V(1,2) < -5.600000E-1)? -6.625000E-3 * V(1,2) - 3.532700E-3:
+ (V(1,2) < -5.400000E-1)? -3.906500E-3 * V(1,2) - 2.010340E-3:
+ (V(1,2) < -5.200000E-1)? -2.222000E-3 * V(1,2) - 1.100710E-3:
+ (V(1,2) < -5.000000E-1)? -1.231000E-3 * V(1,2) - 5.853900E-4:
+ (V(1,2) < -4.800000E-1)? -6.715000E-4 * V(1,2) - 3.056400E-4:
+ (V(1,2) < -4.600000E-1)? -3.660500E-4 * V(1,2) - 1.590240E-4:
+ (V(1,2) < -4.400000E-1)? -2.009000E-4 * V(1,2) - 8.305500E-5:
+ (V(1,2) < -4.200000E-1)? -1.110000E-4 * V(1,2) - 4.349900E-5:
+ (V(1,2) < -4.000000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -3.800000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -3.600000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -3.400000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -3.200000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -3.000000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -2.800000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -2.600000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -2.400000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -2.200000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -2.000000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -1.800000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -1.600000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -1.400000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -1.200000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -1.000000E-1)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -8.000000E-2)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -6.000000E-2)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -4.000000E-2)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < -2.000000E-2)? -0.000000E0 * V(1,2) + 3.121000E-6:
+ (V(1,2) < 0.000000E0)? -1.560500E-4 * V(1,2) + 0.000000E0:
+ 0.000000E0 
.ENDS

* GC BRANCH
.SUBCKT HSTL_II_F_HR_IN50_GND_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -1.500000E0)? -8.430000E-1:
+ (V(1,2) < -1.460000E0)? 1.517500E0 * V(1,2) + 1.433250E0:
+ (V(1,2) < -1.420000E0)? 1.505000E0 * V(1,2) + 1.415000E0:
+ (V(1,2) < -1.380000E0)? 1.492500E0 * V(1,2) + 1.397250E0:
+ (V(1,2) < -1.340000E0)? 1.480000E0 * V(1,2) + 1.380000E0:
+ (V(1,2) < -1.300000E0)? 1.460000E0 * V(1,2) + 1.353200E0:
+ (V(1,2) < -1.260000E0)? 1.435000E0 * V(1,2) + 1.320700E0:
+ (V(1,2) < -1.220000E0)? 1.410000E0 * V(1,2) + 1.289200E0:
+ (V(1,2) < -1.180000E0)? 1.377500E0 * V(1,2) + 1.249550E0:
+ (V(1,2) < -1.140000E0)? 1.337500E0 * V(1,2) + 1.202350E0:
+ (V(1,2) < -1.100000E0)? 1.292500E0 * V(1,2) + 1.151050E0:
+ (V(1,2) < -1.060000E0)? 1.232500E0 * V(1,2) + 1.085050E0:
+ (V(1,2) < -1.020000E0)? 1.140000E0 * V(1,2) + 9.870000E-1:
+ (V(1,2) < -9.800000E-1)? 1.012500E0 * V(1,2) + 8.569500E-1:
+ (V(1,2) < -9.400000E-1)? 8.325000E-1 * V(1,2) + 6.805500E-1:
+ (V(1,2) < -9.000000E-1)? 6.050000E-1 * V(1,2) + 4.667000E-1:
+ (V(1,2) < -8.600000E-1)? 3.892500E-1 * V(1,2) + 2.725250E-1:
+ (V(1,2) < -8.200000E-1)? 2.610000E-1 * V(1,2) + 1.622300E-1:
+ (V(1,2) < -7.800000E-1)? 2.065000E-1 * V(1,2) + 1.175400E-1:
+ (V(1,2) < -7.400000E-1)? 1.832500E-1 * V(1,2) + 9.940500E-2:
+ (V(1,2) < -7.000000E-1)? 1.697500E-1 * V(1,2) + 8.941500E-2:
+ (V(1,2) < -6.600000E-1)? 1.575000E-1 * V(1,2) + 8.084000E-2:
+ (V(1,2) < -6.200000E-1)? 1.437500E-1 * V(1,2) + 7.176500E-2:
+ (V(1,2) < -5.800000E-1)? 1.280000E-1 * V(1,2) + 6.200000E-2:
+ (V(1,2) < -5.400000E-1)? 1.083750E-1 * V(1,2) + 5.061750E-2:
+ (V(1,2) < -5.000000E-1)? 8.490000E-2 * V(1,2) + 3.794100E-2:
+ (V(1,2) < -4.600000E-1)? 5.815000E-2 * V(1,2) + 2.456600E-2:
+ (V(1,2) < -4.200000E-1)? 3.260750E-2 * V(1,2) + 1.281645E-2:
+ (V(1,2) < -3.800000E-1)? 1.445750E-2 * V(1,2) + 5.193450E-3:
+ (V(1,2) < -3.400000E-1)? 5.240000E-3 * V(1,2) + 1.690800E-3:
+ (V(1,2) < -3.000000E-1)? 1.640750E-3 * V(1,2) + 4.670550E-4:
+ (V(1,2) < -2.600000E-1)? 4.644750E-4 * V(1,2) + 1.141725E-4:
+ (V(1,2) < -2.200000E-1)? 1.230250E-4 * V(1,2) + 2.539550E-5:
+ (V(1,2) < -1.800000E-1)? 3.134250E-5 * V(1,2) + 5.225350E-6:
+ (V(1,2) < -1.400000E-1)? 7.802500E-6 * V(1,2) + 9.881500E-7:
+ (V(1,2) < -1.000000E-1)? 1.923500E-6 * V(1,2) + 1.650900E-7:
+ (V(1,2) < -6.000000E-2)? 4.769500E-7 * V(1,2) + 2.043500E-8:
+ (V(1,2) < -2.000000E-2)? 1.256250E-7 * V(1,2) - 6.445000E-10:
+ (V(1,2) < 2.000000E-2)? 3.795000E-8 * V(1,2) - 2.398000E-9:
+ (V(1,2) < 6.000000E-2)? 1.684000E-8 * V(1,2) - 1.975800E-9:
+ (V(1,2) < 1.000000E-1)? 1.032500E-8 * V(1,2) - 1.584900E-9:
+ (V(1,2) < 1.400000E-1)? 8.322500E-9 * V(1,2) - 1.384650E-9:
+ (V(1,2) < 1.800000E-1)? 7.322250E-9 * V(1,2) - 1.244615E-9:
+ (V(1,2) < 2.200000E-1)? 6.497750E-9 * V(1,2) - 1.096205E-9:
+ (V(1,2) < 2.600000E-1)? 6.100000E-9 * V(1,2) - 1.008700E-9:
+ (V(1,2) < 3.000000E-1)? 5.850000E-9 * V(1,2) - 9.437000E-10:
+ (V(1,2) < 3.400000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 3.800000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 4.200000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 4.600000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 5.000000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 5.400000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 5.800000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 6.200000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 6.600000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 7.000000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 7.400000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 7.800000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 8.200000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 8.600000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 9.000000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 9.400000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 9.800000E-1)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.020000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.060000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.100000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.140000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.180000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.220000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.260000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.300000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.340000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.380000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.420000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.460000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ (V(1,2) < 1.500000E0)? -0.000000E0 * V(1,2) + 8.113000E-10:
+ 8.113000E-10 
.ENDS

************************************* END **************************************


.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-0.5

.SUBCKT NOTUSED N1 N2 N3 N4
* NOTHING HERE: OPEN BETWEEN ALL TERMINALS
.ENDS

