

.subckt TL_2 1 2 ngnd length=0.0581254


WTL1 1 ngnd 2 ngnd n=1 RLGCfile=w6l1.rlc l='length'



.ends TL_2
