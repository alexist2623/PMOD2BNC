

.subckt TL_SL2 1 2 ngnd length=0.000127


WTL1 1 ngnd 2 ngnd n=1 RLGCfile=G6Q1.rlc l='length'



.ends TL_SL2
