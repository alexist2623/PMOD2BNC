** Profile: "SCHEMATIC1-Trans"  [ C:\Jeonghyun\GIT\PMOD2BNC\22_1\IBIS_SIM-PSpiceFiles\SCHEMATIC1\Trans.sim ] 

** Creating circuit file "Trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "C:\Jeonghyun\GIT\PMOD2BNC\IBIS\PSPICE\spartan7.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 0.01n 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
