

.subckt R50_withpkg 1 2


R1 1 3 25
R2 3 4 25
Cbody 3 0 1p
Lpkg 4 2 1n


.ends R50_withpkg
