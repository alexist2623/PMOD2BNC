********************************************************************************
*
* LTSPICE MODEL FOR IBIS MODEL(S)
* MODELING DATE: 20230602163639
* GENERAETD BY BPRO: http://www.spisim.com
*
* NOTE: ramp data in .ibs model is used in this converted spice model.
*       VT waveform based conversion will yield more accurate result.
*
********************************************************************************


******************************** BEGIN *****************************************
* ORIG. MDL: C:\Jeonghyun\GIT\PMOD2BNC\IBIS\spartan7_v1.3\spartan7\spartan7.ibs;HSTL_I_F_HR_IN50;TYP
* TERMINALS: INPUT OUTPUT VCC VSS ENABLE

.SUBCKT HSTL_I_F_HR_IN50_TYP NINP NOUT NVCC NVSS NENB

* POWER-ON SOURCE



* INPUT CONTROL
B1 N820 0 V= ((V(NINP) > 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0
B2 N830 0 V= ((V(NINP) < 0.5) & (V(NENB) > 0.5))? 1.0 : 0.0

* RAMP RATE CONTROL
* RISERMP = 4.029756E4 = 0.6318/0.2546n
* FALLRMP = 3.665966E4 = 0.6664/0.2443n

B3 NVCC N850 I= (V(N830) > 0.5)? 0 : V(NVCC, N850) / 3.665966E4
B4 N840 NVSS I= (V(N820) > 0.5)? 0 : V(N840, NVSS) / 4.029756E4
C1 NVCC N850 1F
C2 N840 NVSS 1F
S1 N220 N850 0 N820 SMOD
S2 N840 N220 0 N830 SMOD

G1 N008 NVSS N002 N008 1
G2 NVCC N008 N008 N003 1
R1 N006 NVSS 1
R2 NVCC N006 1

* PU/PD/PC/GC BRANCH
XASRC_PD N002 NVSS N008 N840 HSTL_I_F_HR_IN50_PULLDOWN_TYP
XASRC_PU N003 NVCC N850 N008 HSTL_I_F_HR_IN50_PULLUP_TYP
XASRC_PC N006 NVCC NVCC N006 HSTL_I_F_HR_IN50_POWER_CLAMP_TYP
XASRC_GC N006 NVSS N006 NVSS HSTL_I_F_HR_IN50_GND_CLAMP_TYP

* PACKAGE PARASITICS:
ROPKG N001 NOUT 3.345000E-1
COPKG NOUT NVSS 7.200000E-13
LOPKG N005 N001 4.350000E-9
CCOMP N005 NVSS 7.690000E-12

* Voltage Sources for measuring currents
V5 N006 N005 0
V6 N008 N006 0
V7 N220 N008 0
.ENDS

* PU BRANCH
.SUBCKT HSTL_I_F_HR_IN50_PULLUP_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -1.500000E0)? 4.359500E-2:
+ (V(1,2) < -1.450000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.350000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.250000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.150000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.050000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -9.500000E-1)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -8.500000E-1)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -8.000000E-1)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -7.500000E-1)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -7.000000E-1)? -0.000000E0 * V(1,2) + 4.359500E-2:
+ (V(1,2) < -6.500000E-1)? -4.946000E-2 * V(1,2) + 8.973000E-3:
+ (V(1,2) < -6.000000E-1)? -4.727600E-2 * V(1,2) + 1.039260E-2:
+ (V(1,2) < -5.500000E-1)? -6.467600E-2 * V(1,2) - 4.740000E-5:
+ (V(1,2) < -5.000000E-1)? -6.729800E-2 * V(1,2) - 1.489500E-3:
+ (V(1,2) < -4.500000E-1)? -6.827800E-2 * V(1,2) - 1.979500E-3:
+ (V(1,2) < -4.000000E-1)? -6.785800E-2 * V(1,2) - 1.790500E-3:
+ (V(1,2) < -3.500000E-1)? -6.676200E-2 * V(1,2) - 1.352100E-3:
+ (V(1,2) < -3.000000E-1)? -6.592000E-2 * V(1,2) - 1.057400E-3:
+ (V(1,2) < -2.500000E-1)? -6.477800E-2 * V(1,2) - 7.148000E-4:
+ (V(1,2) < -2.000000E-1)? -6.399600E-2 * V(1,2) - 5.193000E-4:
+ (V(1,2) < -1.500000E-1)? -6.289800E-2 * V(1,2) - 2.997000E-4:
+ (V(1,2) < -1.000000E-1)? -6.210000E-2 * V(1,2) - 1.800000E-4:
+ (V(1,2) < -5.000000E-2)? -6.078000E-2 * V(1,2) - 4.800000E-5:
+ (V(1,2) < 0.000000E0)? -5.845677E-2 * V(1,2) + 6.816140E-5:
+ (V(1,2) < 5.000000E-2)? -5.846323E-2 * V(1,2) + 6.816140E-5:
+ (V(1,2) < 1.000000E-1)? -5.554000E-2 * V(1,2) - 7.800000E-5:
+ (V(1,2) < 1.500000E-1)? -5.074000E-2 * V(1,2) - 5.580000E-4:
+ (V(1,2) < 2.000000E-1)? -4.602000E-2 * V(1,2) - 1.266000E-3:
+ (V(1,2) < 2.500000E-1)? -4.600000E-2 * V(1,2) - 1.270000E-3:
+ (V(1,2) < 3.000000E-1)? -4.600000E-2 * V(1,2) - 1.270000E-3:
+ (V(1,2) < 3.500000E-1)? -4.600000E-2 * V(1,2) - 1.270000E-3:
+ (V(1,2) < 4.000000E-1)? -3.960000E-2 * V(1,2) - 3.510000E-3:
+ (V(1,2) < 4.500000E-1)? -3.640000E-2 * V(1,2) - 4.790000E-3:
+ (V(1,2) < 5.000000E-1)? -3.400000E-2 * V(1,2) - 5.870000E-3:
+ (V(1,2) < 5.500000E-1)? -3.080000E-2 * V(1,2) - 7.470000E-3:
+ (V(1,2) < 6.000000E-1)? -2.720000E-2 * V(1,2) - 9.450000E-3:
+ (V(1,2) < 6.500000E-1)? -2.520000E-2 * V(1,2) - 1.065000E-2:
+ (V(1,2) < 7.000000E-1)? -1.940000E-2 * V(1,2) - 1.442000E-2:
+ (V(1,2) < 7.500000E-1)? -1.920000E-2 * V(1,2) - 1.456000E-2:
+ (V(1,2) < 8.000000E-1)? -1.780000E-2 * V(1,2) - 1.561000E-2:
+ (V(1,2) < 8.500000E-1)? -1.180000E-2 * V(1,2) - 2.041000E-2:
+ (V(1,2) < 9.000000E-1)? -1.200000E-2 * V(1,2) - 2.024000E-2:
+ (V(1,2) < 9.500000E-1)? -1.140000E-2 * V(1,2) - 2.078000E-2:
+ (V(1,2) < 1.000000E0)? -8.000000E-3 * V(1,2) - 2.401000E-2:
+ (V(1,2) < 1.050000E0)? -7.200000E-3 * V(1,2) - 2.481000E-2:
+ (V(1,2) < 1.100000E0)? -6.000000E-3 * V(1,2) - 2.607000E-2:
+ (V(1,2) < 1.150000E0)? -5.400000E-3 * V(1,2) - 2.673000E-2:
+ (V(1,2) < 1.200000E0)? -5.400000E-3 * V(1,2) - 2.673000E-2:
+ (V(1,2) < 1.250000E0)? -4.600000E-3 * V(1,2) - 2.769000E-2:
+ (V(1,2) < 1.300000E0)? -4.400000E-3 * V(1,2) - 2.794000E-2:
+ (V(1,2) < 1.350000E0)? -4.200000E-3 * V(1,2) - 2.820000E-2:
+ (V(1,2) < 1.400000E0)? -4.000000E-3 * V(1,2) - 2.847000E-2:
+ (V(1,2) < 1.450000E0)? -3.600000E-3 * V(1,2) - 2.903000E-2:
+ (V(1,2) < 1.500000E0)? -3.600000E-3 * V(1,2) - 2.903000E-2:
+ (V(1,2) < 1.550000E0)? -3.400000E-3 * V(1,2) - 2.933000E-2:
+ (V(1,2) < 1.600000E0)? -3.200000E-3 * V(1,2) - 2.964000E-2:
+ (V(1,2) < 1.650000E0)? -3.196000E-3 * V(1,2) - 2.964640E-2:
+ (V(1,2) < 1.700000E0)? -3.170000E-3 * V(1,2) - 2.968930E-2:
+ (V(1,2) < 1.750000E0)? -3.140000E-3 * V(1,2) - 2.974030E-2:
+ (V(1,2) < 1.800000E0)? -2.668000E-3 * V(1,2) - 3.056630E-2:
+ (V(1,2) < 1.850000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 1.900000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 1.950000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.000000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.050000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.100000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.150000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.200000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.250000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.300000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.350000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.400000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.450000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.500000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.550000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.600000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.650000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.700000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.750000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.800000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.850000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.900000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 2.950000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ (V(1,2) < 3.000000E0)? -0.000000E0 * V(1,2) - 3.536870E-2:
+ -3.536870E-2
.ENDS

* PD BRANCH
.SUBCKT HSTL_I_F_HR_IN50_PULLDOWN_TYP 3 4 1 2
B1 3 4 V =
+ (V(1,2) < -1.500000E0)? -3.034000E-2:
+ (V(1,2) < -1.450000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.400000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.350000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.300000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.250000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.200000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.150000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.100000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.050000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -1.000000E0)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -9.500000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -9.000000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -8.500000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -8.000000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -7.500000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -7.000000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -6.500000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -6.000000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -5.500000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -5.000000E-1)? -0.000000E0 * V(1,2) - 3.034000E-2:
+ (V(1,2) < -4.500000E-1)? 3.314000E-2 * V(1,2) - 1.377000E-2:
+ (V(1,2) < -4.000000E-1)? 5.448000E-2 * V(1,2) - 4.167000E-3:
+ (V(1,2) < -3.500000E-1)? 5.449000E-2 * V(1,2) - 4.163000E-3:
+ (V(1,2) < -3.000000E-1)? 5.711600E-2 * V(1,2) - 3.243900E-3:
+ (V(1,2) < -2.500000E-1)? 6.326800E-2 * V(1,2) - 1.398300E-3:
+ (V(1,2) < -2.000000E-1)? 6.574000E-2 * V(1,2) - 7.803000E-4:
+ (V(1,2) < -1.500000E-1)? 6.657000E-2 * V(1,2) - 6.143000E-4:
+ (V(1,2) < -1.000000E-1)? 6.871600E-2 * V(1,2) - 2.924000E-4:
+ (V(1,2) < -5.000000E-2)? 7.126000E-2 * V(1,2) - 3.800000E-5:
+ (V(1,2) < 0.000000E0)? 7.184330E-2 * V(1,2) - 8.835100E-6:
+ (V(1,2) < 5.000000E-2)? 7.113670E-2 * V(1,2) - 8.835100E-6:
+ (V(1,2) < 1.000000E-1)? 6.732000E-2 * V(1,2) + 1.820000E-4:
+ (V(1,2) < 1.500000E-1)? 6.232000E-2 * V(1,2) + 6.820000E-4:
+ (V(1,2) < 2.000000E-1)? 5.900000E-2 * V(1,2) + 1.180000E-3:
+ (V(1,2) < 2.500000E-1)? 5.380000E-2 * V(1,2) + 2.220000E-3:
+ (V(1,2) < 3.000000E-1)? 4.920000E-2 * V(1,2) + 3.370000E-3:
+ (V(1,2) < 3.500000E-1)? 4.660000E-2 * V(1,2) + 4.150000E-3:
+ (V(1,2) < 4.000000E-1)? 3.820000E-2 * V(1,2) + 7.090000E-3:
+ (V(1,2) < 4.500000E-1)? 3.820000E-2 * V(1,2) + 7.090000E-3:
+ (V(1,2) < 5.000000E-1)? 3.820000E-2 * V(1,2) + 7.090000E-3:
+ (V(1,2) < 5.500000E-1)? 3.600000E-2 * V(1,2) + 8.190000E-3:
+ (V(1,2) < 6.000000E-1)? 2.820000E-2 * V(1,2) + 1.248000E-2:
+ (V(1,2) < 6.500000E-1)? 2.220000E-2 * V(1,2) + 1.608000E-2:
+ (V(1,2) < 7.000000E-1)? 2.240000E-2 * V(1,2) + 1.595000E-2:
+ (V(1,2) < 7.500000E-1)? 2.020000E-2 * V(1,2) + 1.749000E-2:
+ (V(1,2) < 8.000000E-1)? 1.220000E-2 * V(1,2) + 2.349000E-2:
+ (V(1,2) < 8.500000E-1)? 1.200000E-2 * V(1,2) + 2.365000E-2:
+ (V(1,2) < 9.000000E-1)? 1.220000E-2 * V(1,2) + 2.348000E-2:
+ (V(1,2) < 9.500000E-1)? 1.180000E-2 * V(1,2) + 2.384000E-2:
+ (V(1,2) < 1.000000E0)? 5.000000E-3 * V(1,2) + 3.030000E-2:
+ (V(1,2) < 1.050000E0)? 5.000000E-3 * V(1,2) + 3.030000E-2:
+ (V(1,2) < 1.100000E0)? 5.000000E-3 * V(1,2) + 3.030000E-2:
+ (V(1,2) < 1.150000E0)? 4.800000E-3 * V(1,2) + 3.052000E-2:
+ (V(1,2) < 1.200000E0)? 2.400000E-3 * V(1,2) + 3.328000E-2:
+ (V(1,2) < 1.250000E0)? 1.800000E-3 * V(1,2) + 3.400000E-2:
+ (V(1,2) < 1.300000E0)? 1.200000E-3 * V(1,2) + 3.475000E-2:
+ (V(1,2) < 1.350000E0)? 1.000000E-3 * V(1,2) + 3.501000E-2:
+ (V(1,2) < 1.400000E0)? 1.000000E-3 * V(1,2) + 3.501000E-2:
+ (V(1,2) < 1.450000E0)? 8.000000E-4 * V(1,2) + 3.529000E-2:
+ (V(1,2) < 1.500000E0)? 6.000000E-4 * V(1,2) + 3.558000E-2:
+ (V(1,2) < 1.550000E0)? 6.000000E-4 * V(1,2) + 3.558000E-2:
+ (V(1,2) < 1.600000E0)? 6.000000E-4 * V(1,2) + 3.558000E-2:
+ (V(1,2) < 1.650000E0)? 4.000000E-4 * V(1,2) + 3.590000E-2:
+ (V(1,2) < 1.700000E0)? 3.980000E-4 * V(1,2) + 3.590330E-2:
+ (V(1,2) < 1.750000E0)? 3.940000E-4 * V(1,2) + 3.591010E-2:
+ (V(1,2) < 1.800000E0)? 3.820000E-4 * V(1,2) + 3.593110E-2:
+ (V(1,2) < 1.850000E0)? 3.080000E-4 * V(1,2) + 3.606430E-2:
+ (V(1,2) < 1.900000E0)? 3.660000E-4 * V(1,2) + 3.595700E-2:
+ (V(1,2) < 1.950000E0)? 4.640000E-4 * V(1,2) + 3.577080E-2:
+ (V(1,2) < 2.000000E0)? 6.400000E-5 * V(1,2) + 3.655080E-2:
+ (V(1,2) < 2.050000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.100000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.150000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.200000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.250000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.300000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.350000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.400000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.450000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.500000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.550000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.600000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.650000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.700000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.750000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.800000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.850000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.900000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 2.950000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ (V(1,2) < 3.000000E0)? -0.000000E0 * V(1,2) + 3.667880E-2:
+ 3.667880E-2
.ENDS

* PC BRANCH
.SUBCKT HSTL_I_F_HR_IN50_POWER_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -1.500000E0)? 8.278000E-1:
+ (V(1,2) < -1.480000E0)? -1.535000E0 * V(1,2) - 1.474700E0:
+ (V(1,2) < -1.460000E0)? -1.535000E0 * V(1,2) - 1.474700E0:
+ (V(1,2) < -1.440000E0)? -1.535000E0 * V(1,2) - 1.474700E0:
+ (V(1,2) < -1.420000E0)? -1.530000E0 * V(1,2) - 1.467500E0:
+ (V(1,2) < -1.400000E0)? -1.530000E0 * V(1,2) - 1.467500E0:
+ (V(1,2) < -1.380000E0)? -1.525000E0 * V(1,2) - 1.460500E0:
+ (V(1,2) < -1.360000E0)? -1.530000E0 * V(1,2) - 1.467400E0:
+ (V(1,2) < -1.340000E0)? -1.525000E0 * V(1,2) - 1.460600E0:
+ (V(1,2) < -1.320000E0)? -1.495000E0 * V(1,2) - 1.420400E0:
+ (V(1,2) < -1.300000E0)? -1.500000E0 * V(1,2) - 1.427000E0:
+ (V(1,2) < -1.280000E0)? -1.495000E0 * V(1,2) - 1.420500E0:
+ (V(1,2) < -1.260000E0)? -1.500000E0 * V(1,2) - 1.426900E0:
+ (V(1,2) < -1.240000E0)? -1.490000E0 * V(1,2) - 1.414300E0:
+ (V(1,2) < -1.220000E0)? -1.445000E0 * V(1,2) - 1.358500E0:
+ (V(1,2) < -1.200000E0)? -1.440000E0 * V(1,2) - 1.352400E0:
+ (V(1,2) < -1.180000E0)? -1.445000E0 * V(1,2) - 1.358400E0:
+ (V(1,2) < -1.160000E0)? -1.440000E0 * V(1,2) - 1.352500E0:
+ (V(1,2) < -1.140000E0)? -1.430000E0 * V(1,2) - 1.340900E0:
+ (V(1,2) < -1.120000E0)? -1.325000E0 * V(1,2) - 1.221200E0:
+ (V(1,2) < -1.100000E0)? -1.330000E0 * V(1,2) - 1.226800E0:
+ (V(1,2) < -1.080000E0)? -1.325000E0 * V(1,2) - 1.221300E0:
+ (V(1,2) < -1.060000E0)? -1.325000E0 * V(1,2) - 1.221300E0:
+ (V(1,2) < -1.040000E0)? -1.290000E0 * V(1,2) - 1.184200E0:
+ (V(1,2) < -1.020000E0)? -1.020000E0 * V(1,2) - 9.034000E-1:
+ (V(1,2) < -1.000000E0)? -1.020000E0 * V(1,2) - 9.034000E-1:
+ (V(1,2) < -9.800000E-1)? -1.021000E0 * V(1,2) - 9.044000E-1:
+ (V(1,2) < -9.600000E-1)? -1.020500E0 * V(1,2) - 9.039100E-1:
+ (V(1,2) < -9.400000E-1)? -9.420000E-1 * V(1,2) - 8.285500E-1:
+ (V(1,2) < -9.200000E-1)? -4.085000E-1 * V(1,2) - 3.270600E-1:
+ (V(1,2) < -9.000000E-1)? -4.085000E-1 * V(1,2) - 3.270600E-1:
+ (V(1,2) < -8.800000E-1)? -4.085000E-1 * V(1,2) - 3.270600E-1:
+ (V(1,2) < -8.600000E-1)? -4.090000E-1 * V(1,2) - 3.275000E-1:
+ (V(1,2) < -8.400000E-1)? -3.695000E-1 * V(1,2) - 2.935300E-1:
+ (V(1,2) < -8.200000E-1)? -1.070000E-1 * V(1,2) - 7.303000E-2:
+ (V(1,2) < -8.000000E-1)? -1.065000E-1 * V(1,2) - 7.262000E-2:
+ (V(1,2) < -7.800000E-1)? -1.070000E-1 * V(1,2) - 7.302000E-2:
+ (V(1,2) < -7.600000E-1)? -1.066500E-1 * V(1,2) - 7.274700E-2:
+ (V(1,2) < -7.400000E-1)? -9.950000E-2 * V(1,2) - 6.731300E-2:
+ (V(1,2) < -7.200000E-1)? -5.050000E-2 * V(1,2) - 3.105300E-2:
+ (V(1,2) < -7.000000E-1)? -5.050000E-2 * V(1,2) - 3.105300E-2:
+ (V(1,2) < -6.800000E-1)? -5.045000E-2 * V(1,2) - 3.101800E-2:
+ (V(1,2) < -6.600000E-1)? -5.050000E-2 * V(1,2) - 3.105200E-2:
+ (V(1,2) < -6.400000E-1)? -4.585000E-2 * V(1,2) - 2.798300E-2:
+ (V(1,2) < -6.200000E-1)? -1.435000E-2 * V(1,2) - 7.823000E-3:
+ (V(1,2) < -6.000000E-1)? -1.433000E-2 * V(1,2) - 7.810600E-3:
+ (V(1,2) < -5.800000E-1)? -1.435000E-2 * V(1,2) - 7.822600E-3:
+ (V(1,2) < -5.600000E-1)? -1.434500E-2 * V(1,2) - 7.819700E-3:
+ (V(1,2) < -5.400000E-1)? -4.740000E-3 * V(1,2) - 2.440900E-3:
+ (V(1,2) < -5.200000E-1)? -2.485500E-3 * V(1,2) - 1.223470E-3:
+ (V(1,2) < -5.000000E-1)? -1.853000E-3 * V(1,2) - 8.945700E-4:
+ (V(1,2) < -4.800000E-1)? -7.565000E-4 * V(1,2) - 3.463200E-4:
+ (V(1,2) < -4.600000E-1)? -3.691500E-4 * V(1,2) - 1.603920E-4:
+ (V(1,2) < -4.400000E-1)? -1.947500E-4 * V(1,2) - 8.016800E-5:
+ (V(1,2) < -4.200000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -4.000000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -3.800000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -3.600000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -3.400000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -3.200000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -3.000000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -2.800000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -2.600000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -2.400000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -2.200000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -2.000000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -1.800000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -1.600000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -1.400000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -1.200000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -1.000000E-1)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -8.000000E-2)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -6.000000E-2)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -4.000000E-2)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < -2.000000E-2)? -0.000000E0 * V(1,2) + 5.522000E-6:
+ (V(1,2) < 0.000000E0)? -2.761000E-4 * V(1,2) + 0.000000E0:
+ 0.000000E0
.ENDS

* GC BRANCH
.SUBCKT HSTL_I_F_HR_IN50_GND_CLAMP_TYP 3 4 1 2
B1 3 4 I =
+ (V(1,2) < -1.500000E0)? -8.430000E-1:
+ (V(1,2) < -1.460000E0)? 1.515000E0 * V(1,2) + 1.429500E0:
+ (V(1,2) < -1.420000E0)? 1.500000E0 * V(1,2) + 1.407600E0:
+ (V(1,2) < -1.380000E0)? 1.490000E0 * V(1,2) + 1.393400E0:
+ (V(1,2) < -1.340000E0)? 1.480000E0 * V(1,2) + 1.379600E0:
+ (V(1,2) < -1.300000E0)? 1.410000E0 * V(1,2) + 1.285800E0:
+ (V(1,2) < -1.260000E0)? 1.407500E0 * V(1,2) + 1.282550E0:
+ (V(1,2) < -1.220000E0)? 1.407500E0 * V(1,2) + 1.282550E0:
+ (V(1,2) < -1.180000E0)? 1.410000E0 * V(1,2) + 1.285600E0:
+ (V(1,2) < -1.140000E0)? 1.367500E0 * V(1,2) + 1.235450E0:
+ (V(1,2) < -1.100000E0)? 1.117500E0 * V(1,2) + 9.504500E-1:
+ (V(1,2) < -1.060000E0)? 1.120000E0 * V(1,2) + 9.532000E-1:
+ (V(1,2) < -1.020000E0)? 1.117500E0 * V(1,2) + 9.505500E-1:
+ (V(1,2) < -9.800000E-1)? 1.117500E0 * V(1,2) + 9.505500E-1:
+ (V(1,2) < -9.400000E-1)? 1.047500E0 * V(1,2) + 8.819500E-1:
+ (V(1,2) < -9.000000E-1)? 6.077500E-1 * V(1,2) + 4.685850E-1:
+ (V(1,2) < -8.600000E-1)? 4.005000E-1 * V(1,2) + 2.820600E-1:
+ (V(1,2) < -8.200000E-1)? 2.227500E-1 * V(1,2) + 1.291950E-1:
+ (V(1,2) < -7.800000E-1)? 2.145000E-1 * V(1,2) + 1.224300E-1:
+ (V(1,2) < -7.400000E-1)? 2.145000E-1 * V(1,2) + 1.224300E-1:
+ (V(1,2) < -7.000000E-1)? 1.612500E-1 * V(1,2) + 8.302500E-2:
+ (V(1,2) < -6.600000E-1)? 1.572500E-1 * V(1,2) + 8.022500E-2:
+ (V(1,2) < -6.200000E-1)? 1.505000E-1 * V(1,2) + 7.577000E-2:
+ (V(1,2) < -5.800000E-1)? 9.875000E-2 * V(1,2) + 4.368500E-2:
+ (V(1,2) < -5.400000E-1)? 9.860000E-2 * V(1,2) + 4.359800E-2:
+ (V(1,2) < -5.000000E-1)? 9.870000E-2 * V(1,2) + 4.365200E-2:
+ (V(1,2) < -4.600000E-1)? 8.062500E-2 * V(1,2) + 3.461450E-2:
+ (V(1,2) < -4.200000E-1)? 1.285000E-2 * V(1,2) + 3.438000E-3:
+ (V(1,2) < -3.800000E-1)? 1.287500E-2 * V(1,2) + 3.448500E-3:
+ (V(1,2) < -3.400000E-1)? 1.286000E-2 * V(1,2) + 3.442800E-3:
+ (V(1,2) < -3.000000E-1)? 1.286250E-2 * V(1,2) + 3.443650E-3:
+ (V(1,2) < -2.600000E-1)? 1.018858E-2 * V(1,2) + 2.641473E-3:
+ (V(1,2) < -2.200000E-1)? 1.437250E-4 * V(1,2) + 2.981150E-5:
+ (V(1,2) < -1.800000E-1)? 3.033000E-5 * V(1,2) + 4.864600E-6:
+ (V(1,2) < -1.400000E-1)? 1.155500E-5 * V(1,2) + 1.485100E-6:
+ (V(1,2) < -1.000000E-1)? 2.264250E-6 * V(1,2) + 1.843950E-7:
+ (V(1,2) < -6.000000E-2)? 8.528750E-7 * V(1,2) + 4.325750E-8:
+ (V(1,2) < -2.000000E-2)? 1.221500E-7 * V(1,2) - 5.860000E-10:
+ (V(1,2) < 2.000000E-2)? 3.977500E-8 * V(1,2) - 2.233500E-9:
+ (V(1,2) < 6.000000E-2)? 1.303000E-8 * V(1,2) - 1.698600E-9:
+ (V(1,2) < 1.000000E-1)? 1.302000E-8 * V(1,2) - 1.698000E-9:
+ (V(1,2) < 1.400000E-1)? 1.220675E-8 * V(1,2) - 1.616675E-9:
+ (V(1,2) < 1.800000E-1)? 7.268250E-9 * V(1,2) - 9.252850E-10:
+ (V(1,2) < 2.200000E-1)? 6.592500E-9 * V(1,2) - 8.036500E-10:
+ (V(1,2) < 2.600000E-1)? 6.150000E-9 * V(1,2) - 7.063000E-10:
+ (V(1,2) < 3.000000E-1)? 5.907500E-9 * V(1,2) - 6.432500E-10:
+ (V(1,2) < 3.400000E-1)? 5.525000E-9 * V(1,2) - 5.285000E-10:
+ (V(1,2) < 3.800000E-1)? 5.550000E-9 * V(1,2) - 5.370000E-10:
+ (V(1,2) < 4.200000E-1)? 5.250000E-9 * V(1,2) - 4.230000E-10:
+ (V(1,2) < 4.600000E-1)? 5.050000E-9 * V(1,2) - 3.390000E-10:
+ (V(1,2) < 5.000000E-1)? 5.050000E-9 * V(1,2) - 3.390000E-10:
+ (V(1,2) < 5.400000E-1)? 5.075000E-9 * V(1,2) - 3.515000E-10:
+ (V(1,2) < 5.800000E-1)? 4.925000E-9 * V(1,2) - 2.705000E-10:
+ (V(1,2) < 6.200000E-1)? 4.900000E-9 * V(1,2) - 2.560000E-10:
+ (V(1,2) < 6.600000E-1)? 4.900000E-9 * V(1,2) - 2.560000E-10:
+ (V(1,2) < 7.000000E-1)? 4.900000E-9 * V(1,2) - 2.560000E-10:
+ (V(1,2) < 7.400000E-1)? 4.875000E-9 * V(1,2) - 2.385000E-10:
+ (V(1,2) < 7.800000E-1)? 4.925000E-9 * V(1,2) - 2.755000E-10:
+ (V(1,2) < 8.200000E-1)? 5.025000E-9 * V(1,2) - 3.535000E-10:
+ (V(1,2) < 8.600000E-1)? 4.850000E-9 * V(1,2) - 2.100000E-10:
+ (V(1,2) < 9.000000E-1)? 4.975000E-9 * V(1,2) - 3.175000E-10:
+ (V(1,2) < 9.400000E-1)? 5.175000E-9 * V(1,2) - 4.975000E-10:
+ (V(1,2) < 9.800000E-1)? 5.025000E-9 * V(1,2) - 3.565000E-10:
+ (V(1,2) < 1.020000E0)? 5.100000E-9 * V(1,2) - 4.300000E-10:
+ (V(1,2) < 1.060000E0)? 5.500000E-9 * V(1,2) - 8.380000E-10:
+ (V(1,2) < 1.100000E0)? 5.525000E-9 * V(1,2) - 8.645000E-10:
+ (V(1,2) < 1.140000E0)? 5.500000E-9 * V(1,2) - 8.370000E-10:
+ (V(1,2) < 1.180000E0)? 5.500000E-9 * V(1,2) - 8.370000E-10:
+ (V(1,2) < 1.220000E0)? 6.400000E-9 * V(1,2) - 1.899000E-9:
+ (V(1,2) < 1.260000E0)? 6.650000E-9 * V(1,2) - 2.204000E-9:
+ (V(1,2) < 1.300000E0)? 6.675000E-9 * V(1,2) - 2.235500E-9:
+ (V(1,2) < 1.340000E0)? 6.650000E-9 * V(1,2) - 2.203000E-9:
+ (V(1,2) < 1.380000E0)? 9.900000E-9 * V(1,2) - 6.558000E-9:
+ (V(1,2) < 1.420000E0)? 1.090000E-8 * V(1,2) - 7.938000E-9:
+ (V(1,2) < 1.460000E0)? 1.092500E-8 * V(1,2) - 7.973500E-9:
+ (V(1,2) < 1.500000E0)? 1.092500E-8 * V(1,2) - 7.973500E-9:
+ 8.414000E-9
.ENDS

************************************* END **************************************


.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-0.5

.SUBCKT NOTUSED N1 N2 N3 N4
* NOTHING HERE: OPEN BETWEEN ALL TERMINALS
.ENDS

